-- megafunction wizard: %Pixel Buffer DMA Controller v13.0%
-- GENERATION: XML
-- pixel_buffer_dma_ctrlr.vhd

-- Generated using ACDS version 13.0 156 at 2017.10.30.09:27:42

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pixel_buffer_dma_ctrlr is
	port (
		clk                  : in  std_logic                     := '0';             --             clock_reset.clk
		reset                : in  std_logic                     := '0';             --       clock_reset_reset.reset
		master_readdatavalid : in  std_logic                     := '0';             -- avalon_pixel_dma_master.readdatavalid
		master_waitrequest   : in  std_logic                     := '0';             --                        .waitrequest
		master_address       : out std_logic_vector(31 downto 0);                    --                        .address
		master_arbiterlock   : out std_logic;                                        --                        .lock
		master_read          : out std_logic;                                        --                        .read
		master_readdata      : in  std_logic_vector(7 downto 0)  := (others => '0'); --                        .readdata
		slave_address        : in  std_logic_vector(1 downto 0)  := (others => '0'); --    avalon_control_slave.address
		slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => '0'); --                        .byteenable
		slave_read           : in  std_logic                     := '0';             --                        .read
		slave_write          : in  std_logic                     := '0';             --                        .write
		slave_writedata      : in  std_logic_vector(31 downto 0) := (others => '0'); --                        .writedata
		slave_readdata       : out std_logic_vector(31 downto 0);                    --                        .readdata
		stream_ready         : in  std_logic                     := '0';             --     avalon_pixel_source.ready
		stream_startofpacket : out std_logic;                                        --                        .startofpacket
		stream_endofpacket   : out std_logic;                                        --                        .endofpacket
		stream_valid         : out std_logic;                                        --                        .valid
		stream_data          : out std_logic_vector(7 downto 0)                      --                        .data
	);
end entity pixel_buffer_dma_ctrlr;

architecture rtl of pixel_buffer_dma_ctrlr is
	component pixel_buffer_dma_ctrlr_0002 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component pixel_buffer_dma_ctrlr_0002;

begin

	pixel_buffer_dma_ctrlr_inst : component pixel_buffer_dma_ctrlr_0002
		port map (
			clk                  => clk,                  --             clock_reset.clk
			reset                => reset,                --       clock_reset_reset.reset
			master_readdatavalid => master_readdatavalid, -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => master_waitrequest,   --                        .waitrequest
			master_address       => master_address,       --                        .address
			master_arbiterlock   => master_arbiterlock,   --                        .lock
			master_read          => master_read,          --                        .read
			master_readdata      => master_readdata,      --                        .readdata
			slave_address        => slave_address,        --    avalon_control_slave.address
			slave_byteenable     => slave_byteenable,     --                        .byteenable
			slave_read           => slave_read,           --                        .read
			slave_write          => slave_write,          --                        .write
			slave_writedata      => slave_writedata,      --                        .writedata
			slave_readdata       => slave_readdata,       --                        .readdata
			stream_ready         => stream_ready,         --     avalon_pixel_source.ready
			stream_startofpacket => stream_startofpacket, --                        .startofpacket
			stream_endofpacket   => stream_endofpacket,   --                        .endofpacket
			stream_valid         => stream_valid,         --                        .valid
			stream_data          => stream_data           --                        .data
		);

end architecture rtl; -- of pixel_buffer_dma_ctrlr
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2017 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_up_avalon_video_pixel_buffer_dma" version="13.0" >
-- Retrieval info: 	<generic name="addr_mode" value="X-Y" />
-- Retrieval info: 	<generic name="start_address" value="0" />
-- Retrieval info: 	<generic name="back_start_address" value="0" />
-- Retrieval info: 	<generic name="image_width" value="640" />
-- Retrieval info: 	<generic name="image_height" value="480" />
-- Retrieval info: 	<generic name="color_space" value="8-bit Grayscale" />
-- Retrieval info: 	<generic name="AUTO_CLOCK_RESET_CLOCK_RATE" value="-1" />
-- Retrieval info: 	<generic name="AUTO_DEVICE_FAMILY" value="Cyclone IV GX" />
-- Retrieval info: </instance>
-- IPFS_FILES : pixel_buffer_dma_ctrlr.vho
-- RELATED_FILES: pixel_buffer_dma_ctrlr.vhd, pixel_buffer_dma_ctrlr_0002.v
