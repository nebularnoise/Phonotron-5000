-- nios_ii.vhd

-- Generated using ACDS version 13.0 156 at 2017.11.13.16:17:28

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nios_ii is
	port (
		sram_de2_ADDR            : out   std_logic_vector(17 downto 0);                    --       sram_de2.ADDR
		sram_de2_DQ              : inout std_logic_vector(15 downto 0) := (others => '0'); --               .DQ
		sram_de2_WE_N            : out   std_logic;                                        --               .WE_N
		sram_de2_OE_N            : out   std_logic;                                        --               .OE_N
		sram_de2_UB_N            : out   std_logic;                                        --               .UB_N
		sram_de2_LB_N            : out   std_logic;                                        --               .LB_N
		sram_de2_CE_N            : out   std_logic;                                        --               .CE_N
		color_out_export         : out   std_logic_vector(1 downto 0);                     --      color_out.export
		wr_address_export        : out   std_logic_vector(16 downto 0);                    --     wr_address.export
		seq_clap_export          : out   std_logic_vector(31 downto 0);                    --       seq_clap.export
		seq_kick_export          : out   std_logic_vector(31 downto 0);                    --       seq_kick.export
		wr_en_export             : out   std_logic;                                        --          wr_en.export
		reset_100_reset_n        : in    std_logic                     := '0';             --      reset_100.reset_n
		in_bus_export            : in    std_logic_vector(19 downto 0) := (others => '0'); --         in_bus.export
		clk_100_clk              : in    std_logic                     := '0';             --        clk_100.clk
		led_r_export             : out   std_logic_vector(17 downto 0);                    --          led_r.export
		seq_snare_export         : out   std_logic_vector(31 downto 0);                    --      seq_snare.export
		seq_hh_export            : out   std_logic_vector(31 downto 0);                    --         seq_hh.export
		kb_data_export           : in    std_logic_vector(7 downto 0)  := (others => '0'); --        kb_data.export
		kb_irq_export            : in    std_logic                     := '0';             --         kb_irq.export
		kick_irq_export          : in    std_logic                     := '0';             --       kick_irq.export
		snare_irq_export         : in    std_logic                     := '0';             --      snare_irq.export
		hh_irq_export            : in    std_logic                     := '0';             --         hh_irq.export
		clap_irq_export          : in    std_logic                     := '0';             --       clap_irq.export
		dac_irq_export           : in    std_logic                     := '0';             --        dac_irq.export
		audio_dac_fifo_oAUD_BCK  : out   std_logic;                                        -- audio_dac_fifo.oAUD_BCK
		audio_dac_fifo_oAUD_LRCK : out   std_logic;                                        --               .oAUD_LRCK
		audio_dac_fifo_oAUD_DATA : out   std_logic;                                        --               .oAUD_DATA
		audio_dac_fifo_oAUD_XCK  : out   std_logic;                                        --               .oAUD_XCK
		audio_dac_fifo_iCLK_18_4 : in    std_logic                     := '0';             --               .iCLK_18_4
		audio_sos_export         : out   std_logic_vector(31 downto 0)                     --      audio_sos.export
	);
end entity nios_ii;

architecture rtl of nios_ii is
	component SRAM_DE2 is
		port (
			clk               : in    std_logic                     := 'X';             -- clk
			reset_n           : in    std_logic                     := 'X';             -- reset_n
			avs_s0_readdata   : out   std_logic_vector(15 downto 0);                    -- readdata
			avs_s0_writedata  : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avs_s0_address    : in    std_logic_vector(17 downto 0) := (others => 'X'); -- address
			avs_s0_write      : in    std_logic                     := 'X';             -- write
			avs_s0_read       : in    std_logic                     := 'X';             -- read
			avs_s0_byteenable : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			coe_SRAM_ADDR     : out   std_logic_vector(17 downto 0);                    -- export
			coe_SRAM_DQ       : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			coe_SRAM_WE_N     : out   std_logic;                                        -- export
			coe_SRAM_OE_N     : out   std_logic;                                        -- export
			coe_SRAM_UB_N     : out   std_logic;                                        -- export
			coe_SRAM_LB_N     : out   std_logic;                                        -- export
			coe_SRAM_CE_N     : out   std_logic                                         -- export
		);
	end component SRAM_DE2;

	component nios_ii_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(20 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(20 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component nios_ii_nios2_qsys_0;

	component nios_ii_in_bus is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(19 downto 0) := (others => 'X')  -- export
		);
	end component nios_ii_in_bus;

	component nios_ii_wr_en is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component nios_ii_wr_en;

	component nios_ii_color_out is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component nios_ii_color_out;

	component nios_ii_wr_address is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(16 downto 0)                     -- export
		);
	end component nios_ii_wr_address;

	component nios_ii_seq_clap is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component nios_ii_seq_clap;

	component nios_ii_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component nios_ii_timer_0;

	component nios_ii_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component nios_ii_jtag_uart_0;

	component nios_ii_led_r is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component nios_ii_led_r;

	component nios_ii_kb_irq is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component nios_ii_kb_irq;

	component nios_ii_kb_data is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component nios_ii_kb_data;

	component AUDIO_DAC_FIFO is
		generic (
			REF_CLK     : integer := 18432000;
			SAMPLE_RATE : integer := 8000;
			DATA_WIDTH  : integer := 16;
			CHANNEL_NUM : integer := 2
		);
		port (
			avs_s0_writedata : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avs_s0_write     : in  std_logic                     := 'X';             -- write
			avs_s0_readdata  : out std_logic_vector(15 downto 0);                    -- readdata
			avs_s0_read      : in  std_logic                     := 'X';             -- read
			clk              : in  std_logic                     := 'X';             -- clk
			reset_n          : in  std_logic                     := 'X';             -- reset_n
			oAUD_BCK         : out std_logic;                                        -- export
			oAUD_LRCK        : out std_logic;                                        -- export
			oAUD_DATA        : out std_logic;                                        -- export
			oAUD_XCK         : out std_logic;                                        -- export
			iCLK_18_4        : in  std_logic                     := 'X'              -- export
		);
	end component AUDIO_DAC_FIFO;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(97 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component nios_ii_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(97 downto 0);                    -- data
			src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_ii_addr_router;

	component nios_ii_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(97 downto 0);                    -- data
			src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_ii_addr_router_001;

	component nios_ii_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(97 downto 0);                    -- data
			src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_ii_id_router;

	component nios_ii_id_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(79 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(79 downto 0);                    -- data
			src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_ii_id_router_001;

	component nios_ii_id_router_020 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(97 downto 0);                    -- data
			src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_ii_id_router_020;

	component nios_ii_id_router_021 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(79 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(79 downto 0);                    -- data
			src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component nios_ii_id_router_021;

	component altera_merlin_traffic_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                        -- ready
			cmd_sink_valid         : in  std_logic                     := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                     := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(97 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			cmd_src_startofpacket  : out std_logic;                                        -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                        -- endofpacket
			rsp_sink_ready         : out std_logic;                                        -- ready
			rsp_sink_valid         : in  std_logic                     := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                     := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                        -- valid
			rsp_src_data           : out std_logic_vector(97 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(22 downto 0);                    -- channel
			rsp_src_startofpacket  : out std_logic;                                        -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                        -- endofpacket
			cmd_src_valid          : out std_logic_vector(22 downto 0)                     -- data
		);
	end component altera_merlin_traffic_limiter;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(79 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(79 downto 0);                    -- data
			source0_channel       : out std_logic_vector(22 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component nios_ii_cmd_xbar_demux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			sink_ready          : out std_logic;                                        -- ready
			sink_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(22 downto 0) := (others => 'X'); -- data
			src0_ready          : in  std_logic                     := 'X';             -- ready
			src0_valid          : out std_logic;                                        -- valid
			src0_data           : out std_logic_vector(97 downto 0);                    -- data
			src0_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src0_startofpacket  : out std_logic;                                        -- startofpacket
			src0_endofpacket    : out std_logic;                                        -- endofpacket
			src1_ready          : in  std_logic                     := 'X';             -- ready
			src1_valid          : out std_logic;                                        -- valid
			src1_data           : out std_logic_vector(97 downto 0);                    -- data
			src1_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src1_startofpacket  : out std_logic;                                        -- startofpacket
			src1_endofpacket    : out std_logic;                                        -- endofpacket
			src2_ready          : in  std_logic                     := 'X';             -- ready
			src2_valid          : out std_logic;                                        -- valid
			src2_data           : out std_logic_vector(97 downto 0);                    -- data
			src2_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src2_startofpacket  : out std_logic;                                        -- startofpacket
			src2_endofpacket    : out std_logic;                                        -- endofpacket
			src3_ready          : in  std_logic                     := 'X';             -- ready
			src3_valid          : out std_logic;                                        -- valid
			src3_data           : out std_logic_vector(97 downto 0);                    -- data
			src3_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src3_startofpacket  : out std_logic;                                        -- startofpacket
			src3_endofpacket    : out std_logic;                                        -- endofpacket
			src4_ready          : in  std_logic                     := 'X';             -- ready
			src4_valid          : out std_logic;                                        -- valid
			src4_data           : out std_logic_vector(97 downto 0);                    -- data
			src4_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src4_startofpacket  : out std_logic;                                        -- startofpacket
			src4_endofpacket    : out std_logic;                                        -- endofpacket
			src5_ready          : in  std_logic                     := 'X';             -- ready
			src5_valid          : out std_logic;                                        -- valid
			src5_data           : out std_logic_vector(97 downto 0);                    -- data
			src5_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src5_startofpacket  : out std_logic;                                        -- startofpacket
			src5_endofpacket    : out std_logic;                                        -- endofpacket
			src6_ready          : in  std_logic                     := 'X';             -- ready
			src6_valid          : out std_logic;                                        -- valid
			src6_data           : out std_logic_vector(97 downto 0);                    -- data
			src6_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src6_startofpacket  : out std_logic;                                        -- startofpacket
			src6_endofpacket    : out std_logic;                                        -- endofpacket
			src7_ready          : in  std_logic                     := 'X';             -- ready
			src7_valid          : out std_logic;                                        -- valid
			src7_data           : out std_logic_vector(97 downto 0);                    -- data
			src7_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src7_startofpacket  : out std_logic;                                        -- startofpacket
			src7_endofpacket    : out std_logic;                                        -- endofpacket
			src8_ready          : in  std_logic                     := 'X';             -- ready
			src8_valid          : out std_logic;                                        -- valid
			src8_data           : out std_logic_vector(97 downto 0);                    -- data
			src8_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src8_startofpacket  : out std_logic;                                        -- startofpacket
			src8_endofpacket    : out std_logic;                                        -- endofpacket
			src9_ready          : in  std_logic                     := 'X';             -- ready
			src9_valid          : out std_logic;                                        -- valid
			src9_data           : out std_logic_vector(97 downto 0);                    -- data
			src9_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src9_startofpacket  : out std_logic;                                        -- startofpacket
			src9_endofpacket    : out std_logic;                                        -- endofpacket
			src10_ready         : in  std_logic                     := 'X';             -- ready
			src10_valid         : out std_logic;                                        -- valid
			src10_data          : out std_logic_vector(97 downto 0);                    -- data
			src10_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src10_startofpacket : out std_logic;                                        -- startofpacket
			src10_endofpacket   : out std_logic;                                        -- endofpacket
			src11_ready         : in  std_logic                     := 'X';             -- ready
			src11_valid         : out std_logic;                                        -- valid
			src11_data          : out std_logic_vector(97 downto 0);                    -- data
			src11_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src11_startofpacket : out std_logic;                                        -- startofpacket
			src11_endofpacket   : out std_logic;                                        -- endofpacket
			src12_ready         : in  std_logic                     := 'X';             -- ready
			src12_valid         : out std_logic;                                        -- valid
			src12_data          : out std_logic_vector(97 downto 0);                    -- data
			src12_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src12_startofpacket : out std_logic;                                        -- startofpacket
			src12_endofpacket   : out std_logic;                                        -- endofpacket
			src13_ready         : in  std_logic                     := 'X';             -- ready
			src13_valid         : out std_logic;                                        -- valid
			src13_data          : out std_logic_vector(97 downto 0);                    -- data
			src13_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src13_startofpacket : out std_logic;                                        -- startofpacket
			src13_endofpacket   : out std_logic;                                        -- endofpacket
			src14_ready         : in  std_logic                     := 'X';             -- ready
			src14_valid         : out std_logic;                                        -- valid
			src14_data          : out std_logic_vector(97 downto 0);                    -- data
			src14_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src14_startofpacket : out std_logic;                                        -- startofpacket
			src14_endofpacket   : out std_logic;                                        -- endofpacket
			src15_ready         : in  std_logic                     := 'X';             -- ready
			src15_valid         : out std_logic;                                        -- valid
			src15_data          : out std_logic_vector(97 downto 0);                    -- data
			src15_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src15_startofpacket : out std_logic;                                        -- startofpacket
			src15_endofpacket   : out std_logic;                                        -- endofpacket
			src16_ready         : in  std_logic                     := 'X';             -- ready
			src16_valid         : out std_logic;                                        -- valid
			src16_data          : out std_logic_vector(97 downto 0);                    -- data
			src16_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src16_startofpacket : out std_logic;                                        -- startofpacket
			src16_endofpacket   : out std_logic;                                        -- endofpacket
			src17_ready         : in  std_logic                     := 'X';             -- ready
			src17_valid         : out std_logic;                                        -- valid
			src17_data          : out std_logic_vector(97 downto 0);                    -- data
			src17_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src17_startofpacket : out std_logic;                                        -- startofpacket
			src17_endofpacket   : out std_logic;                                        -- endofpacket
			src18_ready         : in  std_logic                     := 'X';             -- ready
			src18_valid         : out std_logic;                                        -- valid
			src18_data          : out std_logic_vector(97 downto 0);                    -- data
			src18_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src18_startofpacket : out std_logic;                                        -- startofpacket
			src18_endofpacket   : out std_logic;                                        -- endofpacket
			src19_ready         : in  std_logic                     := 'X';             -- ready
			src19_valid         : out std_logic;                                        -- valid
			src19_data          : out std_logic_vector(97 downto 0);                    -- data
			src19_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src19_startofpacket : out std_logic;                                        -- startofpacket
			src19_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios_ii_cmd_xbar_demux;

	component nios_ii_cmd_xbar_demux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			sink_ready          : out std_logic;                                        -- ready
			sink_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(22 downto 0) := (others => 'X'); -- data
			src0_ready          : in  std_logic                     := 'X';             -- ready
			src0_valid          : out std_logic;                                        -- valid
			src0_data           : out std_logic_vector(97 downto 0);                    -- data
			src0_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src0_startofpacket  : out std_logic;                                        -- startofpacket
			src0_endofpacket    : out std_logic;                                        -- endofpacket
			src1_ready          : in  std_logic                     := 'X';             -- ready
			src1_valid          : out std_logic;                                        -- valid
			src1_data           : out std_logic_vector(97 downto 0);                    -- data
			src1_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src1_startofpacket  : out std_logic;                                        -- startofpacket
			src1_endofpacket    : out std_logic;                                        -- endofpacket
			src2_ready          : in  std_logic                     := 'X';             -- ready
			src2_valid          : out std_logic;                                        -- valid
			src2_data           : out std_logic_vector(97 downto 0);                    -- data
			src2_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src2_startofpacket  : out std_logic;                                        -- startofpacket
			src2_endofpacket    : out std_logic;                                        -- endofpacket
			src3_ready          : in  std_logic                     := 'X';             -- ready
			src3_valid          : out std_logic;                                        -- valid
			src3_data           : out std_logic_vector(97 downto 0);                    -- data
			src3_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src3_startofpacket  : out std_logic;                                        -- startofpacket
			src3_endofpacket    : out std_logic;                                        -- endofpacket
			src4_ready          : in  std_logic                     := 'X';             -- ready
			src4_valid          : out std_logic;                                        -- valid
			src4_data           : out std_logic_vector(97 downto 0);                    -- data
			src4_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src4_startofpacket  : out std_logic;                                        -- startofpacket
			src4_endofpacket    : out std_logic;                                        -- endofpacket
			src5_ready          : in  std_logic                     := 'X';             -- ready
			src5_valid          : out std_logic;                                        -- valid
			src5_data           : out std_logic_vector(97 downto 0);                    -- data
			src5_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src5_startofpacket  : out std_logic;                                        -- startofpacket
			src5_endofpacket    : out std_logic;                                        -- endofpacket
			src6_ready          : in  std_logic                     := 'X';             -- ready
			src6_valid          : out std_logic;                                        -- valid
			src6_data           : out std_logic_vector(97 downto 0);                    -- data
			src6_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src6_startofpacket  : out std_logic;                                        -- startofpacket
			src6_endofpacket    : out std_logic;                                        -- endofpacket
			src7_ready          : in  std_logic                     := 'X';             -- ready
			src7_valid          : out std_logic;                                        -- valid
			src7_data           : out std_logic_vector(97 downto 0);                    -- data
			src7_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src7_startofpacket  : out std_logic;                                        -- startofpacket
			src7_endofpacket    : out std_logic;                                        -- endofpacket
			src8_ready          : in  std_logic                     := 'X';             -- ready
			src8_valid          : out std_logic;                                        -- valid
			src8_data           : out std_logic_vector(97 downto 0);                    -- data
			src8_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src8_startofpacket  : out std_logic;                                        -- startofpacket
			src8_endofpacket    : out std_logic;                                        -- endofpacket
			src9_ready          : in  std_logic                     := 'X';             -- ready
			src9_valid          : out std_logic;                                        -- valid
			src9_data           : out std_logic_vector(97 downto 0);                    -- data
			src9_channel        : out std_logic_vector(22 downto 0);                    -- channel
			src9_startofpacket  : out std_logic;                                        -- startofpacket
			src9_endofpacket    : out std_logic;                                        -- endofpacket
			src10_ready         : in  std_logic                     := 'X';             -- ready
			src10_valid         : out std_logic;                                        -- valid
			src10_data          : out std_logic_vector(97 downto 0);                    -- data
			src10_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src10_startofpacket : out std_logic;                                        -- startofpacket
			src10_endofpacket   : out std_logic;                                        -- endofpacket
			src11_ready         : in  std_logic                     := 'X';             -- ready
			src11_valid         : out std_logic;                                        -- valid
			src11_data          : out std_logic_vector(97 downto 0);                    -- data
			src11_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src11_startofpacket : out std_logic;                                        -- startofpacket
			src11_endofpacket   : out std_logic;                                        -- endofpacket
			src12_ready         : in  std_logic                     := 'X';             -- ready
			src12_valid         : out std_logic;                                        -- valid
			src12_data          : out std_logic_vector(97 downto 0);                    -- data
			src12_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src12_startofpacket : out std_logic;                                        -- startofpacket
			src12_endofpacket   : out std_logic;                                        -- endofpacket
			src13_ready         : in  std_logic                     := 'X';             -- ready
			src13_valid         : out std_logic;                                        -- valid
			src13_data          : out std_logic_vector(97 downto 0);                    -- data
			src13_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src13_startofpacket : out std_logic;                                        -- startofpacket
			src13_endofpacket   : out std_logic;                                        -- endofpacket
			src14_ready         : in  std_logic                     := 'X';             -- ready
			src14_valid         : out std_logic;                                        -- valid
			src14_data          : out std_logic_vector(97 downto 0);                    -- data
			src14_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src14_startofpacket : out std_logic;                                        -- startofpacket
			src14_endofpacket   : out std_logic;                                        -- endofpacket
			src15_ready         : in  std_logic                     := 'X';             -- ready
			src15_valid         : out std_logic;                                        -- valid
			src15_data          : out std_logic_vector(97 downto 0);                    -- data
			src15_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src15_startofpacket : out std_logic;                                        -- startofpacket
			src15_endofpacket   : out std_logic;                                        -- endofpacket
			src16_ready         : in  std_logic                     := 'X';             -- ready
			src16_valid         : out std_logic;                                        -- valid
			src16_data          : out std_logic_vector(97 downto 0);                    -- data
			src16_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src16_startofpacket : out std_logic;                                        -- startofpacket
			src16_endofpacket   : out std_logic;                                        -- endofpacket
			src17_ready         : in  std_logic                     := 'X';             -- ready
			src17_valid         : out std_logic;                                        -- valid
			src17_data          : out std_logic_vector(97 downto 0);                    -- data
			src17_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src17_startofpacket : out std_logic;                                        -- startofpacket
			src17_endofpacket   : out std_logic;                                        -- endofpacket
			src18_ready         : in  std_logic                     := 'X';             -- ready
			src18_valid         : out std_logic;                                        -- valid
			src18_data          : out std_logic_vector(97 downto 0);                    -- data
			src18_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src18_startofpacket : out std_logic;                                        -- startofpacket
			src18_endofpacket   : out std_logic;                                        -- endofpacket
			src19_ready         : in  std_logic                     := 'X';             -- ready
			src19_valid         : out std_logic;                                        -- valid
			src19_data          : out std_logic_vector(97 downto 0);                    -- data
			src19_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src19_startofpacket : out std_logic;                                        -- startofpacket
			src19_endofpacket   : out std_logic;                                        -- endofpacket
			src20_ready         : in  std_logic                     := 'X';             -- ready
			src20_valid         : out std_logic;                                        -- valid
			src20_data          : out std_logic_vector(97 downto 0);                    -- data
			src20_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src20_startofpacket : out std_logic;                                        -- startofpacket
			src20_endofpacket   : out std_logic;                                        -- endofpacket
			src21_ready         : in  std_logic                     := 'X';             -- ready
			src21_valid         : out std_logic;                                        -- valid
			src21_data          : out std_logic_vector(97 downto 0);                    -- data
			src21_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src21_startofpacket : out std_logic;                                        -- startofpacket
			src21_endofpacket   : out std_logic;                                        -- endofpacket
			src22_ready         : in  std_logic                     := 'X';             -- ready
			src22_valid         : out std_logic;                                        -- valid
			src22_data          : out std_logic_vector(97 downto 0);                    -- data
			src22_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src22_startofpacket : out std_logic;                                        -- startofpacket
			src22_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios_ii_cmd_xbar_demux_001;

	component nios_ii_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(97 downto 0);                    -- data
			src_channel         : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios_ii_cmd_xbar_mux;

	component nios_ii_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(97 downto 0);                    -- data
			src0_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(97 downto 0);                    -- data
			src1_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios_ii_rsp_xbar_demux;

	component nios_ii_rsp_xbar_demux_020 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(97 downto 0);                    -- data
			src0_channel       : out std_logic_vector(22 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component nios_ii_rsp_xbar_demux_020;

	component nios_ii_rsp_xbar_mux is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			src_ready            : in  std_logic                     := 'X';             -- ready
			src_valid            : out std_logic;                                        -- valid
			src_data             : out std_logic_vector(97 downto 0);                    -- data
			src_channel          : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket    : out std_logic;                                        -- startofpacket
			src_endofpacket      : out std_logic;                                        -- endofpacket
			sink0_ready          : out std_logic;                                        -- ready
			sink0_valid          : in  std_logic                     := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                        -- ready
			sink1_valid          : in  std_logic                     := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                        -- ready
			sink2_valid          : in  std_logic                     := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                        -- ready
			sink3_valid          : in  std_logic                     := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                        -- ready
			sink4_valid          : in  std_logic                     := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                        -- ready
			sink5_valid          : in  std_logic                     := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                        -- ready
			sink6_valid          : in  std_logic                     := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                        -- ready
			sink7_valid          : in  std_logic                     := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                        -- ready
			sink8_valid          : in  std_logic                     := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                        -- ready
			sink9_valid          : in  std_logic                     := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                        -- ready
			sink10_valid         : in  std_logic                     := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                        -- ready
			sink11_valid         : in  std_logic                     := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                        -- ready
			sink12_valid         : in  std_logic                     := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                        -- ready
			sink13_valid         : in  std_logic                     := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink14_ready         : out std_logic;                                        -- ready
			sink14_valid         : in  std_logic                     := 'X';             -- valid
			sink14_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink14_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink14_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink14_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink15_ready         : out std_logic;                                        -- ready
			sink15_valid         : in  std_logic                     := 'X';             -- valid
			sink15_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink15_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink15_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink15_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink16_ready         : out std_logic;                                        -- ready
			sink16_valid         : in  std_logic                     := 'X';             -- valid
			sink16_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink16_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink16_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink16_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink17_ready         : out std_logic;                                        -- ready
			sink17_valid         : in  std_logic                     := 'X';             -- valid
			sink17_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink17_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink17_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink17_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink18_ready         : out std_logic;                                        -- ready
			sink18_valid         : in  std_logic                     := 'X';             -- valid
			sink18_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink18_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink18_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink18_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink19_ready         : out std_logic;                                        -- ready
			sink19_valid         : in  std_logic                     := 'X';             -- valid
			sink19_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink19_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink19_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink19_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios_ii_rsp_xbar_mux;

	component nios_ii_rsp_xbar_mux_001 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			src_ready            : in  std_logic                     := 'X';             -- ready
			src_valid            : out std_logic;                                        -- valid
			src_data             : out std_logic_vector(97 downto 0);                    -- data
			src_channel          : out std_logic_vector(22 downto 0);                    -- channel
			src_startofpacket    : out std_logic;                                        -- startofpacket
			src_endofpacket      : out std_logic;                                        -- endofpacket
			sink0_ready          : out std_logic;                                        -- ready
			sink0_valid          : in  std_logic                     := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                        -- ready
			sink1_valid          : in  std_logic                     := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                        -- ready
			sink2_valid          : in  std_logic                     := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                        -- ready
			sink3_valid          : in  std_logic                     := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                        -- ready
			sink4_valid          : in  std_logic                     := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                        -- ready
			sink5_valid          : in  std_logic                     := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                        -- ready
			sink6_valid          : in  std_logic                     := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                        -- ready
			sink7_valid          : in  std_logic                     := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                        -- ready
			sink8_valid          : in  std_logic                     := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                        -- ready
			sink9_valid          : in  std_logic                     := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                        -- ready
			sink10_valid         : in  std_logic                     := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                        -- ready
			sink11_valid         : in  std_logic                     := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                        -- ready
			sink12_valid         : in  std_logic                     := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                        -- ready
			sink13_valid         : in  std_logic                     := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink14_ready         : out std_logic;                                        -- ready
			sink14_valid         : in  std_logic                     := 'X';             -- valid
			sink14_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink14_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink14_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink14_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink15_ready         : out std_logic;                                        -- ready
			sink15_valid         : in  std_logic                     := 'X';             -- valid
			sink15_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink15_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink15_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink15_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink16_ready         : out std_logic;                                        -- ready
			sink16_valid         : in  std_logic                     := 'X';             -- valid
			sink16_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink16_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink16_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink16_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink17_ready         : out std_logic;                                        -- ready
			sink17_valid         : in  std_logic                     := 'X';             -- valid
			sink17_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink17_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink17_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink17_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink18_ready         : out std_logic;                                        -- ready
			sink18_valid         : in  std_logic                     := 'X';             -- valid
			sink18_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink18_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink18_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink18_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink19_ready         : out std_logic;                                        -- ready
			sink19_valid         : in  std_logic                     := 'X';             -- valid
			sink19_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink19_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink19_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink19_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink20_ready         : out std_logic;                                        -- ready
			sink20_valid         : in  std_logic                     := 'X';             -- valid
			sink20_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink20_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink20_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink20_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink21_ready         : out std_logic;                                        -- ready
			sink21_valid         : in  std_logic                     := 'X';             -- valid
			sink21_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink21_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink21_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink21_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink22_ready         : out std_logic;                                        -- ready
			sink22_valid         : in  std_logic                     := 'X';             -- valid
			sink22_channel       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			sink22_data          : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			sink22_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink22_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component nios_ii_rsp_xbar_mux_001;

	component nios_ii_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			receiver8_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component nios_ii_irq_mapper;

	component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(98 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(80 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(80 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(20 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(97 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(98 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(20 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(79 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(79 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(80 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(80 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent;

	component nios_ii_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(97 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(79 downto 0);                    -- data
			out_channel          : out std_logic_vector(22 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component nios_ii_width_adapter;

	component nios_ii_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(22 downto 0) := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(79 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(97 downto 0);                    -- data
			out_channel          : out std_logic_vector(22 downto 0);                    -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component nios_ii_width_adapter_001;

	component nios_ii_nios2_qsys_0_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(20 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios_ii_nios2_qsys_0_instruction_master_translator;

	component nios_ii_nios2_qsys_0_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(20 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component nios_ii_nios2_qsys_0_data_master_translator;

	component nios_ii_nios2_qsys_0_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_nios2_qsys_0_jtag_debug_module_translator;

	component nios_ii_sram_de2_0_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(17 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_sram_de2_0_s0_translator;

	component nios_ii_jtag_uart_0_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_jtag_uart_0_avalon_jtag_slave_translator;

	component nios_ii_audio_sos_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_audio_sos_s1_translator;

	component nios_ii_timer_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_timer_0_s1_translator;

	component nios_ii_in_bus_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_in_bus_s1_translator;

	component nios_ii_audio_dac_fifo_0_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component nios_ii_audio_dac_fifo_0_s0_translator;

	signal nios2_qsys_0_instruction_master_waitrequest                                                         : std_logic;                     -- nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                                                             : std_logic_vector(20 downto 0); -- nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	signal nios2_qsys_0_instruction_master_read                                                                : std_logic;                     -- nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	signal nios2_qsys_0_instruction_master_readdata                                                            : std_logic_vector(31 downto 0); -- nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_instruction_master_readdatavalid                                                       : std_logic;                     -- nios2_qsys_0_instruction_master_translator:av_readdatavalid -> nios2_qsys_0:i_readdatavalid
	signal nios2_qsys_0_data_master_waitrequest                                                                : std_logic;                     -- nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_writedata                                                                  : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	signal nios2_qsys_0_data_master_address                                                                    : std_logic_vector(20 downto 0); -- nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	signal nios2_qsys_0_data_master_write                                                                      : std_logic;                     -- nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	signal nios2_qsys_0_data_master_read                                                                       : std_logic;                     -- nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	signal nios2_qsys_0_data_master_readdata                                                                   : std_logic_vector(31 downto 0); -- nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_debugaccess                                                                : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	signal nios2_qsys_0_data_master_readdatavalid                                                              : std_logic;                     -- nios2_qsys_0_data_master_translator:av_readdatavalid -> nios2_qsys_0:d_readdatavalid
	signal nios2_qsys_0_data_master_byteenable                                                                 : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address                               : std_logic_vector(8 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read                                  : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal sram_de2_0_s0_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(15 downto 0); -- SRAM_DE2_0_s0_translator:av_writedata -> SRAM_DE2_0:avs_s0_writedata
	signal sram_de2_0_s0_translator_avalon_anti_slave_0_address                                                : std_logic_vector(17 downto 0); -- SRAM_DE2_0_s0_translator:av_address -> SRAM_DE2_0:avs_s0_address
	signal sram_de2_0_s0_translator_avalon_anti_slave_0_write                                                  : std_logic;                     -- SRAM_DE2_0_s0_translator:av_write -> SRAM_DE2_0:avs_s0_write
	signal sram_de2_0_s0_translator_avalon_anti_slave_0_read                                                   : std_logic;                     -- SRAM_DE2_0_s0_translator:av_read -> SRAM_DE2_0:avs_s0_read
	signal sram_de2_0_s0_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(15 downto 0); -- SRAM_DE2_0:avs_s0_readdata -> SRAM_DE2_0_s0_translator:av_readdata
	signal sram_de2_0_s0_translator_avalon_anti_slave_0_byteenable                                             : std_logic_vector(1 downto 0);  -- SRAM_DE2_0_s0_translator:av_byteenable -> SRAM_DE2_0:avs_s0_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                            : std_logic;                     -- jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(31 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                : std_logic_vector(0 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                             : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                  : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                   : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	signal audio_sos_s1_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(31 downto 0); -- audio_sos_s1_translator:av_writedata -> audio_sos:writedata
	signal audio_sos_s1_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(1 downto 0);  -- audio_sos_s1_translator:av_address -> audio_sos:address
	signal audio_sos_s1_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                     -- audio_sos_s1_translator:av_chipselect -> audio_sos:chipselect
	signal audio_sos_s1_translator_avalon_anti_slave_0_write                                                   : std_logic;                     -- audio_sos_s1_translator:av_write -> audio_sos_s1_translator_avalon_anti_slave_0_write:in
	signal audio_sos_s1_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0); -- audio_sos:readdata -> audio_sos_s1_translator:av_readdata
	signal dac_irq_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0); -- dac_irq_s1_translator:av_writedata -> dac_irq:writedata
	signal dac_irq_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);  -- dac_irq_s1_translator:av_address -> dac_irq:address
	signal dac_irq_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                     -- dac_irq_s1_translator:av_chipselect -> dac_irq:chipselect
	signal dac_irq_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                     -- dac_irq_s1_translator:av_write -> dac_irq_s1_translator_avalon_anti_slave_0_write:in
	signal dac_irq_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0); -- dac_irq:readdata -> dac_irq_s1_translator:av_readdata
	signal clap_irq_s1_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(31 downto 0); -- clap_irq_s1_translator:av_writedata -> clap_irq:writedata
	signal clap_irq_s1_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(1 downto 0);  -- clap_irq_s1_translator:av_address -> clap_irq:address
	signal clap_irq_s1_translator_avalon_anti_slave_0_chipselect                                               : std_logic;                     -- clap_irq_s1_translator:av_chipselect -> clap_irq:chipselect
	signal clap_irq_s1_translator_avalon_anti_slave_0_write                                                    : std_logic;                     -- clap_irq_s1_translator:av_write -> clap_irq_s1_translator_avalon_anti_slave_0_write:in
	signal clap_irq_s1_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0); -- clap_irq:readdata -> clap_irq_s1_translator:av_readdata
	signal hh_irq_s1_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(31 downto 0); -- hh_irq_s1_translator:av_writedata -> hh_irq:writedata
	signal hh_irq_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);  -- hh_irq_s1_translator:av_address -> hh_irq:address
	signal hh_irq_s1_translator_avalon_anti_slave_0_chipselect                                                 : std_logic;                     -- hh_irq_s1_translator:av_chipselect -> hh_irq:chipselect
	signal hh_irq_s1_translator_avalon_anti_slave_0_write                                                      : std_logic;                     -- hh_irq_s1_translator:av_write -> hh_irq_s1_translator_avalon_anti_slave_0_write:in
	signal hh_irq_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0); -- hh_irq:readdata -> hh_irq_s1_translator:av_readdata
	signal snare_irq_s1_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(31 downto 0); -- snare_irq_s1_translator:av_writedata -> snare_irq:writedata
	signal snare_irq_s1_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(1 downto 0);  -- snare_irq_s1_translator:av_address -> snare_irq:address
	signal snare_irq_s1_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                     -- snare_irq_s1_translator:av_chipselect -> snare_irq:chipselect
	signal snare_irq_s1_translator_avalon_anti_slave_0_write                                                   : std_logic;                     -- snare_irq_s1_translator:av_write -> snare_irq_s1_translator_avalon_anti_slave_0_write:in
	signal snare_irq_s1_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0); -- snare_irq:readdata -> snare_irq_s1_translator:av_readdata
	signal kick_irq_s1_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(31 downto 0); -- kick_irq_s1_translator:av_writedata -> kick_irq:writedata
	signal kick_irq_s1_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(1 downto 0);  -- kick_irq_s1_translator:av_address -> kick_irq:address
	signal kick_irq_s1_translator_avalon_anti_slave_0_chipselect                                               : std_logic;                     -- kick_irq_s1_translator:av_chipselect -> kick_irq:chipselect
	signal kick_irq_s1_translator_avalon_anti_slave_0_write                                                    : std_logic;                     -- kick_irq_s1_translator:av_write -> kick_irq_s1_translator_avalon_anti_slave_0_write:in
	signal kick_irq_s1_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0); -- kick_irq:readdata -> kick_irq_s1_translator:av_readdata
	signal kb_irq_s1_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(31 downto 0); -- kb_irq_s1_translator:av_writedata -> kb_irq:writedata
	signal kb_irq_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);  -- kb_irq_s1_translator:av_address -> kb_irq:address
	signal kb_irq_s1_translator_avalon_anti_slave_0_chipselect                                                 : std_logic;                     -- kb_irq_s1_translator:av_chipselect -> kb_irq:chipselect
	signal kb_irq_s1_translator_avalon_anti_slave_0_write                                                      : std_logic;                     -- kb_irq_s1_translator:av_write -> kb_irq_s1_translator_avalon_anti_slave_0_write:in
	signal kb_irq_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0); -- kb_irq:readdata -> kb_irq_s1_translator:av_readdata
	signal seq_hh_s1_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(31 downto 0); -- seq_hh_s1_translator:av_writedata -> seq_hh:writedata
	signal seq_hh_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);  -- seq_hh_s1_translator:av_address -> seq_hh:address
	signal seq_hh_s1_translator_avalon_anti_slave_0_chipselect                                                 : std_logic;                     -- seq_hh_s1_translator:av_chipselect -> seq_hh:chipselect
	signal seq_hh_s1_translator_avalon_anti_slave_0_write                                                      : std_logic;                     -- seq_hh_s1_translator:av_write -> seq_hh_s1_translator_avalon_anti_slave_0_write:in
	signal seq_hh_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0); -- seq_hh:readdata -> seq_hh_s1_translator:av_readdata
	signal seq_snare_s1_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(31 downto 0); -- seq_snare_s1_translator:av_writedata -> seq_snare:writedata
	signal seq_snare_s1_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(1 downto 0);  -- seq_snare_s1_translator:av_address -> seq_snare:address
	signal seq_snare_s1_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                     -- seq_snare_s1_translator:av_chipselect -> seq_snare:chipselect
	signal seq_snare_s1_translator_avalon_anti_slave_0_write                                                   : std_logic;                     -- seq_snare_s1_translator:av_write -> seq_snare_s1_translator_avalon_anti_slave_0_write:in
	signal seq_snare_s1_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0); -- seq_snare:readdata -> seq_snare_s1_translator:av_readdata
	signal led_r_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0); -- led_r_s1_translator:av_writedata -> led_r:writedata
	signal led_r_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);  -- led_r_s1_translator:av_address -> led_r:address
	signal led_r_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                     -- led_r_s1_translator:av_chipselect -> led_r:chipselect
	signal led_r_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                     -- led_r_s1_translator:av_write -> led_r_s1_translator_avalon_anti_slave_0_write:in
	signal led_r_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0); -- led_r:readdata -> led_r_s1_translator:av_readdata
	signal timer_0_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(15 downto 0); -- timer_0_s1_translator:av_writedata -> timer_0:writedata
	signal timer_0_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(2 downto 0);  -- timer_0_s1_translator:av_address -> timer_0:address
	signal timer_0_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                     -- timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	signal timer_0_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                     -- timer_0_s1_translator:av_write -> timer_0_s1_translator_avalon_anti_slave_0_write:in
	signal timer_0_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(15 downto 0); -- timer_0:readdata -> timer_0_s1_translator:av_readdata
	signal seq_clap_s1_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(31 downto 0); -- seq_clap_s1_translator:av_writedata -> seq_clap:writedata
	signal seq_clap_s1_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(1 downto 0);  -- seq_clap_s1_translator:av_address -> seq_clap:address
	signal seq_clap_s1_translator_avalon_anti_slave_0_chipselect                                               : std_logic;                     -- seq_clap_s1_translator:av_chipselect -> seq_clap:chipselect
	signal seq_clap_s1_translator_avalon_anti_slave_0_write                                                    : std_logic;                     -- seq_clap_s1_translator:av_write -> seq_clap_s1_translator_avalon_anti_slave_0_write:in
	signal seq_clap_s1_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0); -- seq_clap:readdata -> seq_clap_s1_translator:av_readdata
	signal seq_kick_s1_translator_avalon_anti_slave_0_writedata                                                : std_logic_vector(31 downto 0); -- seq_kick_s1_translator:av_writedata -> seq_kick:writedata
	signal seq_kick_s1_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(1 downto 0);  -- seq_kick_s1_translator:av_address -> seq_kick:address
	signal seq_kick_s1_translator_avalon_anti_slave_0_chipselect                                               : std_logic;                     -- seq_kick_s1_translator:av_chipselect -> seq_kick:chipselect
	signal seq_kick_s1_translator_avalon_anti_slave_0_write                                                    : std_logic;                     -- seq_kick_s1_translator:av_write -> seq_kick_s1_translator_avalon_anti_slave_0_write:in
	signal seq_kick_s1_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0); -- seq_kick:readdata -> seq_kick_s1_translator:av_readdata
	signal wr_address_s1_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(31 downto 0); -- wr_address_s1_translator:av_writedata -> wr_address:writedata
	signal wr_address_s1_translator_avalon_anti_slave_0_address                                                : std_logic_vector(1 downto 0);  -- wr_address_s1_translator:av_address -> wr_address:address
	signal wr_address_s1_translator_avalon_anti_slave_0_chipselect                                             : std_logic;                     -- wr_address_s1_translator:av_chipselect -> wr_address:chipselect
	signal wr_address_s1_translator_avalon_anti_slave_0_write                                                  : std_logic;                     -- wr_address_s1_translator:av_write -> wr_address_s1_translator_avalon_anti_slave_0_write:in
	signal wr_address_s1_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(31 downto 0); -- wr_address:readdata -> wr_address_s1_translator:av_readdata
	signal color_out_s1_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(31 downto 0); -- color_out_s1_translator:av_writedata -> color_out:writedata
	signal color_out_s1_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(1 downto 0);  -- color_out_s1_translator:av_address -> color_out:address
	signal color_out_s1_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                     -- color_out_s1_translator:av_chipselect -> color_out:chipselect
	signal color_out_s1_translator_avalon_anti_slave_0_write                                                   : std_logic;                     -- color_out_s1_translator:av_write -> color_out_s1_translator_avalon_anti_slave_0_write:in
	signal color_out_s1_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0); -- color_out:readdata -> color_out_s1_translator:av_readdata
	signal in_bus_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);  -- in_bus_s1_translator:av_address -> in_bus:address
	signal in_bus_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0); -- in_bus:readdata -> in_bus_s1_translator:av_readdata
	signal wr_en_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0); -- wr_en_s1_translator:av_writedata -> wr_en:writedata
	signal wr_en_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);  -- wr_en_s1_translator:av_address -> wr_en:address
	signal wr_en_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                     -- wr_en_s1_translator:av_chipselect -> wr_en:chipselect
	signal wr_en_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                     -- wr_en_s1_translator:av_write -> wr_en_s1_translator_avalon_anti_slave_0_write:in
	signal wr_en_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0); -- wr_en:readdata -> wr_en_s1_translator:av_readdata
	signal kb_data_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);  -- kb_data_s1_translator:av_address -> kb_data:address
	signal kb_data_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0); -- kb_data:readdata -> kb_data_s1_translator:av_readdata
	signal audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(15 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator:av_writedata -> AUDIO_DAC_FIFO_0:avs_s0_writedata
	signal audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_write                                            : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator:av_write -> AUDIO_DAC_FIFO_0:avs_s0_write
	signal audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_read                                             : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator:av_read -> AUDIO_DAC_FIFO_0:avs_s0_read
	signal audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(15 downto 0); -- AUDIO_DAC_FIFO_0:avs_s0_readdata -> AUDIO_DAC_FIFO_0_s0_translator:av_readdata
	signal timer_1_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(15 downto 0); -- timer_1_s1_translator:av_writedata -> timer_1:writedata
	signal timer_1_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(2 downto 0);  -- timer_1_s1_translator:av_address -> timer_1:address
	signal timer_1_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                     -- timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	signal timer_1_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                     -- timer_1_s1_translator:av_write -> timer_1_s1_translator_avalon_anti_slave_0_write:in
	signal timer_1_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(15 downto 0); -- timer_1:readdata -> timer_1_s1_translator:av_readdata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest                    : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount                     : std_logic_vector(2 downto 0);  -- nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata                      : std_logic_vector(31 downto 0); -- nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address                        : std_logic_vector(20 downto 0); -- nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock                           : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write                          : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read                           : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata                       : std_logic_vector(31 downto 0); -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess                    : std_logic;                     -- nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable                     : std_logic_vector(3 downto 0);  -- nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid                  : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest                           : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount                            : std_logic_vector(2 downto 0);  -- nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata                             : std_logic_vector(31 downto 0); -- nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_address                               : std_logic_vector(20 downto 0); -- nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock                                  : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_write                                 : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_read                                  : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata                              : std_logic_vector(31 downto 0); -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess                           : std_logic;                     -- nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable                            : std_logic_vector(3 downto 0);  -- nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid                         : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(20 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(98 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(98 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                     -- SRAM_DE2_0_s0_translator:uav_waitrequest -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(1 downto 0);  -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> SRAM_DE2_0_s0_translator:uav_burstcount
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(15 downto 0); -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> SRAM_DE2_0_s0_translator:uav_writedata
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(20 downto 0); -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> SRAM_DE2_0_s0_translator:uav_address
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> SRAM_DE2_0_s0_translator:uav_write
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> SRAM_DE2_0_s0_translator:uav_lock
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> SRAM_DE2_0_s0_translator:uav_read
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(15 downto 0); -- SRAM_DE2_0_s0_translator:uav_readdata -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                     -- SRAM_DE2_0_s0_translator:uav_readdatavalid -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SRAM_DE2_0_s0_translator:uav_debugaccess
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(1 downto 0);  -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> SRAM_DE2_0_s0_translator:uav_byteenable
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(80 downto 0); -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(80 downto 0); -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(17 downto 0); -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(2 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(31 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(20 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(31 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(3 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(98 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(98 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(33 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                     -- audio_sos_s1_translator:uav_waitrequest -> audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);  -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> audio_sos_s1_translator:uav_burstcount
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0); -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> audio_sos_s1_translator:uav_writedata
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(20 downto 0); -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_address -> audio_sos_s1_translator:uav_address
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_write -> audio_sos_s1_translator:uav_write
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_lock -> audio_sos_s1_translator:uav_lock
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_read -> audio_sos_s1_translator:uav_read
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0); -- audio_sos_s1_translator:uav_readdata -> audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                     -- audio_sos_s1_translator:uav_readdatavalid -> audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> audio_sos_s1_translator:uav_debugaccess
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);  -- audio_sos_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> audio_sos_s1_translator:uav_byteenable
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(98 downto 0); -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(98 downto 0); -- audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0); -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                     -- dac_irq_s1_translator:uav_waitrequest -> dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);  -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> dac_irq_s1_translator:uav_burstcount
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0); -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> dac_irq_s1_translator:uav_writedata
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(20 downto 0); -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_address -> dac_irq_s1_translator:uav_address
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_write -> dac_irq_s1_translator:uav_write
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> dac_irq_s1_translator:uav_lock
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_read -> dac_irq_s1_translator:uav_read
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0); -- dac_irq_s1_translator:uav_readdata -> dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                     -- dac_irq_s1_translator:uav_readdatavalid -> dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dac_irq_s1_translator:uav_debugaccess
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);  -- dac_irq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> dac_irq_s1_translator:uav_byteenable
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(98 downto 0); -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(98 downto 0); -- dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0); -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                     -- clap_irq_s1_translator:uav_waitrequest -> clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);  -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> clap_irq_s1_translator:uav_burstcount
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0); -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> clap_irq_s1_translator:uav_writedata
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(20 downto 0); -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_address -> clap_irq_s1_translator:uav_address
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_write -> clap_irq_s1_translator:uav_write
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> clap_irq_s1_translator:uav_lock
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_read -> clap_irq_s1_translator:uav_read
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0); -- clap_irq_s1_translator:uav_readdata -> clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                     -- clap_irq_s1_translator:uav_readdatavalid -> clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> clap_irq_s1_translator:uav_debugaccess
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);  -- clap_irq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> clap_irq_s1_translator:uav_byteenable
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(98 downto 0); -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(98 downto 0); -- clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0); -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                     -- hh_irq_s1_translator:uav_waitrequest -> hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);  -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hh_irq_s1_translator:uav_burstcount
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0); -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hh_irq_s1_translator:uav_writedata
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(20 downto 0); -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_address -> hh_irq_s1_translator:uav_address
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_write -> hh_irq_s1_translator:uav_write
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hh_irq_s1_translator:uav_lock
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_read -> hh_irq_s1_translator:uav_read
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0); -- hh_irq_s1_translator:uav_readdata -> hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                     -- hh_irq_s1_translator:uav_readdatavalid -> hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hh_irq_s1_translator:uav_debugaccess
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- hh_irq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hh_irq_s1_translator:uav_byteenable
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(98 downto 0); -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(98 downto 0); -- hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0); -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                     -- snare_irq_s1_translator:uav_waitrequest -> snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);  -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> snare_irq_s1_translator:uav_burstcount
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0); -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> snare_irq_s1_translator:uav_writedata
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(20 downto 0); -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_address -> snare_irq_s1_translator:uav_address
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_write -> snare_irq_s1_translator:uav_write
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> snare_irq_s1_translator:uav_lock
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_read -> snare_irq_s1_translator:uav_read
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0); -- snare_irq_s1_translator:uav_readdata -> snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                     -- snare_irq_s1_translator:uav_readdatavalid -> snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> snare_irq_s1_translator:uav_debugaccess
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);  -- snare_irq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> snare_irq_s1_translator:uav_byteenable
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(98 downto 0); -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(98 downto 0); -- snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0); -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                     -- kick_irq_s1_translator:uav_waitrequest -> kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);  -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> kick_irq_s1_translator:uav_burstcount
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0); -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> kick_irq_s1_translator:uav_writedata
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(20 downto 0); -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_address -> kick_irq_s1_translator:uav_address
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_write -> kick_irq_s1_translator:uav_write
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> kick_irq_s1_translator:uav_lock
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_read -> kick_irq_s1_translator:uav_read
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0); -- kick_irq_s1_translator:uav_readdata -> kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                     -- kick_irq_s1_translator:uav_readdatavalid -> kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> kick_irq_s1_translator:uav_debugaccess
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);  -- kick_irq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> kick_irq_s1_translator:uav_byteenable
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(98 downto 0); -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(98 downto 0); -- kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0); -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                     -- kb_irq_s1_translator:uav_waitrequest -> kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);  -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> kb_irq_s1_translator:uav_burstcount
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0); -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> kb_irq_s1_translator:uav_writedata
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(20 downto 0); -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_address -> kb_irq_s1_translator:uav_address
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_write -> kb_irq_s1_translator:uav_write
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_lock -> kb_irq_s1_translator:uav_lock
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_read -> kb_irq_s1_translator:uav_read
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0); -- kb_irq_s1_translator:uav_readdata -> kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                     -- kb_irq_s1_translator:uav_readdatavalid -> kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> kb_irq_s1_translator:uav_debugaccess
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- kb_irq_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> kb_irq_s1_translator:uav_byteenable
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(98 downto 0); -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(98 downto 0); -- kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0); -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                     -- seq_hh_s1_translator:uav_waitrequest -> seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);  -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> seq_hh_s1_translator:uav_burstcount
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0); -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> seq_hh_s1_translator:uav_writedata
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(20 downto 0); -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_address -> seq_hh_s1_translator:uav_address
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_write -> seq_hh_s1_translator:uav_write
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_lock -> seq_hh_s1_translator:uav_lock
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_read -> seq_hh_s1_translator:uav_read
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0); -- seq_hh_s1_translator:uav_readdata -> seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                     -- seq_hh_s1_translator:uav_readdatavalid -> seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seq_hh_s1_translator:uav_debugaccess
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- seq_hh_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> seq_hh_s1_translator:uav_byteenable
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(98 downto 0); -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(98 downto 0); -- seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0); -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                     -- seq_snare_s1_translator:uav_waitrequest -> seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);  -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> seq_snare_s1_translator:uav_burstcount
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0); -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> seq_snare_s1_translator:uav_writedata
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(20 downto 0); -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_address -> seq_snare_s1_translator:uav_address
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_write -> seq_snare_s1_translator:uav_write
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_lock -> seq_snare_s1_translator:uav_lock
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_read -> seq_snare_s1_translator:uav_read
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0); -- seq_snare_s1_translator:uav_readdata -> seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                     -- seq_snare_s1_translator:uav_readdatavalid -> seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seq_snare_s1_translator:uav_debugaccess
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);  -- seq_snare_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> seq_snare_s1_translator:uav_byteenable
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(98 downto 0); -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(98 downto 0); -- seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0); -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                     -- led_r_s1_translator:uav_waitrequest -> led_r_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);  -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_r_s1_translator:uav_burstcount
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0); -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_r_s1_translator:uav_writedata
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(20 downto 0); -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_r_s1_translator:uav_address
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_r_s1_translator:uav_write
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_r_s1_translator:uav_lock
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_r_s1_translator:uav_read
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0); -- led_r_s1_translator:uav_readdata -> led_r_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                     -- led_r_s1_translator:uav_readdatavalid -> led_r_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_r_s1_translator:uav_debugaccess
	signal led_r_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);  -- led_r_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_r_s1_translator:uav_byteenable
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(98 downto 0); -- led_r_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_r_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_r_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_r_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_r_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(98 downto 0); -- led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_r_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_r_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0); -- led_r_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_r_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_r_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                     -- timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(20 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0); -- timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                     -- timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(98 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(98 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                     -- seq_clap_s1_translator:uav_waitrequest -> seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);  -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> seq_clap_s1_translator:uav_burstcount
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0); -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> seq_clap_s1_translator:uav_writedata
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(20 downto 0); -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_address -> seq_clap_s1_translator:uav_address
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_write -> seq_clap_s1_translator:uav_write
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_lock -> seq_clap_s1_translator:uav_lock
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_read -> seq_clap_s1_translator:uav_read
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0); -- seq_clap_s1_translator:uav_readdata -> seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                     -- seq_clap_s1_translator:uav_readdatavalid -> seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seq_clap_s1_translator:uav_debugaccess
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);  -- seq_clap_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> seq_clap_s1_translator:uav_byteenable
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(98 downto 0); -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(98 downto 0); -- seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0); -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                     -- seq_kick_s1_translator:uav_waitrequest -> seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);  -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> seq_kick_s1_translator:uav_burstcount
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0); -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> seq_kick_s1_translator:uav_writedata
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(20 downto 0); -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_address -> seq_kick_s1_translator:uav_address
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_write -> seq_kick_s1_translator:uav_write
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_lock -> seq_kick_s1_translator:uav_lock
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_read -> seq_kick_s1_translator:uav_read
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0); -- seq_kick_s1_translator:uav_readdata -> seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                     -- seq_kick_s1_translator:uav_readdatavalid -> seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seq_kick_s1_translator:uav_debugaccess
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);  -- seq_kick_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> seq_kick_s1_translator:uav_byteenable
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(98 downto 0); -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(98 downto 0); -- seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(33 downto 0); -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                     -- wr_address_s1_translator:uav_waitrequest -> wr_address_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);  -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> wr_address_s1_translator:uav_burstcount
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0); -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> wr_address_s1_translator:uav_writedata
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(20 downto 0); -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_address -> wr_address_s1_translator:uav_address
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_write -> wr_address_s1_translator:uav_write
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_lock -> wr_address_s1_translator:uav_lock
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_read -> wr_address_s1_translator:uav_read
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0); -- wr_address_s1_translator:uav_readdata -> wr_address_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                     -- wr_address_s1_translator:uav_readdatavalid -> wr_address_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> wr_address_s1_translator:uav_debugaccess
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);  -- wr_address_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> wr_address_s1_translator:uav_byteenable
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(98 downto 0); -- wr_address_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> wr_address_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> wr_address_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> wr_address_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> wr_address_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(98 downto 0); -- wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> wr_address_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> wr_address_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(33 downto 0); -- wr_address_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> wr_address_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> wr_address_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                     -- color_out_s1_translator:uav_waitrequest -> color_out_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);  -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> color_out_s1_translator:uav_burstcount
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0); -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> color_out_s1_translator:uav_writedata
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(20 downto 0); -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_address -> color_out_s1_translator:uav_address
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_write -> color_out_s1_translator:uav_write
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_lock -> color_out_s1_translator:uav_lock
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_read -> color_out_s1_translator:uav_read
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0); -- color_out_s1_translator:uav_readdata -> color_out_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                     -- color_out_s1_translator:uav_readdatavalid -> color_out_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> color_out_s1_translator:uav_debugaccess
	signal color_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);  -- color_out_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> color_out_s1_translator:uav_byteenable
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(98 downto 0); -- color_out_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> color_out_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> color_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> color_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> color_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(98 downto 0); -- color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> color_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> color_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0); -- color_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> color_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> color_out_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                     -- in_bus_s1_translator:uav_waitrequest -> in_bus_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);  -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> in_bus_s1_translator:uav_burstcount
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0); -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> in_bus_s1_translator:uav_writedata
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(20 downto 0); -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_address -> in_bus_s1_translator:uav_address
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_write -> in_bus_s1_translator:uav_write
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_lock -> in_bus_s1_translator:uav_lock
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_read -> in_bus_s1_translator:uav_read
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0); -- in_bus_s1_translator:uav_readdata -> in_bus_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                     -- in_bus_s1_translator:uav_readdatavalid -> in_bus_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> in_bus_s1_translator:uav_debugaccess
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- in_bus_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> in_bus_s1_translator:uav_byteenable
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(98 downto 0); -- in_bus_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> in_bus_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> in_bus_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> in_bus_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> in_bus_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(98 downto 0); -- in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> in_bus_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> in_bus_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0); -- in_bus_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> in_bus_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> in_bus_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                     -- wr_en_s1_translator:uav_waitrequest -> wr_en_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);  -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> wr_en_s1_translator:uav_burstcount
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0); -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> wr_en_s1_translator:uav_writedata
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(20 downto 0); -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_address -> wr_en_s1_translator:uav_address
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_write -> wr_en_s1_translator:uav_write
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_lock -> wr_en_s1_translator:uav_lock
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_read -> wr_en_s1_translator:uav_read
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0); -- wr_en_s1_translator:uav_readdata -> wr_en_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                     -- wr_en_s1_translator:uav_readdatavalid -> wr_en_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> wr_en_s1_translator:uav_debugaccess
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);  -- wr_en_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> wr_en_s1_translator:uav_byteenable
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(98 downto 0); -- wr_en_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> wr_en_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> wr_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> wr_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> wr_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(98 downto 0); -- wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> wr_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> wr_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0); -- wr_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> wr_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> wr_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                     -- kb_data_s1_translator:uav_waitrequest -> kb_data_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);  -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> kb_data_s1_translator:uav_burstcount
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0); -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> kb_data_s1_translator:uav_writedata
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(20 downto 0); -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_address -> kb_data_s1_translator:uav_address
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_write -> kb_data_s1_translator:uav_write
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_lock -> kb_data_s1_translator:uav_lock
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_read -> kb_data_s1_translator:uav_read
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0); -- kb_data_s1_translator:uav_readdata -> kb_data_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                     -- kb_data_s1_translator:uav_readdatavalid -> kb_data_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> kb_data_s1_translator:uav_debugaccess
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);  -- kb_data_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> kb_data_s1_translator:uav_byteenable
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(98 downto 0); -- kb_data_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> kb_data_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> kb_data_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> kb_data_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> kb_data_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(98 downto 0); -- kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> kb_data_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> kb_data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0); -- kb_data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> kb_data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> kb_data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator:uav_waitrequest -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(1 downto 0);  -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> AUDIO_DAC_FIFO_0_s0_translator:uav_burstcount
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(15 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> AUDIO_DAC_FIFO_0_s0_translator:uav_writedata
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(20 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> AUDIO_DAC_FIFO_0_s0_translator:uav_address
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> AUDIO_DAC_FIFO_0_s0_translator:uav_write
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> AUDIO_DAC_FIFO_0_s0_translator:uav_lock
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> AUDIO_DAC_FIFO_0_s0_translator:uav_read
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(15 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator:uav_readdata -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator:uav_readdatavalid -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> AUDIO_DAC_FIFO_0_s0_translator:uav_debugaccess
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(1 downto 0);  -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> AUDIO_DAC_FIFO_0_s0_translator:uav_byteenable
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(80 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(80 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(17 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                     -- timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(20 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0); -- timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                     -- timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(98 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(98 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket           : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                 : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket         : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data                  : std_logic_vector(97 downto 0); -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                 : std_logic;                     -- addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                  : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid                        : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data                         : std_logic_vector(97 downto 0); -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready                        : std_logic;                     -- addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(97 downto 0); -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(79 downto 0); -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                     -- id_router_001:sink_ready -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(97 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                     -- id_router_002:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(97 downto 0); -- audio_sos_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                     -- id_router_003:sink_ready -> audio_sos_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(97 downto 0); -- dac_irq_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                     -- id_router_004:sink_ready -> dac_irq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(97 downto 0); -- clap_irq_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                     -- id_router_005:sink_ready -> clap_irq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(97 downto 0); -- hh_irq_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                     -- id_router_006:sink_ready -> hh_irq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(97 downto 0); -- snare_irq_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                     -- id_router_007:sink_ready -> snare_irq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(97 downto 0); -- kick_irq_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                     -- id_router_008:sink_ready -> kick_irq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(97 downto 0); -- kb_irq_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                     -- id_router_009:sink_ready -> kb_irq_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(97 downto 0); -- seq_hh_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                     -- id_router_010:sink_ready -> seq_hh_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(97 downto 0); -- seq_snare_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                     -- id_router_011:sink_ready -> seq_snare_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(97 downto 0); -- led_r_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal led_r_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                     -- id_router_012:sink_ready -> led_r_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(97 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                     -- id_router_013:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(97 downto 0); -- seq_clap_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                     -- id_router_014:sink_ready -> seq_clap_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(97 downto 0); -- seq_kick_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	signal seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                     -- id_router_015:sink_ready -> seq_kick_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(97 downto 0); -- wr_address_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	signal wr_address_s1_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                     -- id_router_016:sink_ready -> wr_address_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(97 downto 0); -- color_out_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	signal color_out_s1_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                     -- id_router_017:sink_ready -> color_out_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(97 downto 0); -- in_bus_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	signal in_bus_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                     -- id_router_018:sink_ready -> in_bus_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(97 downto 0); -- wr_en_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	signal wr_en_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                     -- id_router_019:sink_ready -> wr_en_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(97 downto 0); -- kb_data_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	signal kb_data_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                     -- id_router_020:sink_ready -> kb_data_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(79 downto 0); -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	signal audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                     -- id_router_021:sink_ready -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(97 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                     -- id_router_022:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                         : std_logic;                     -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                               : std_logic;                     -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                       : std_logic;                     -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                                : std_logic_vector(97 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                             : std_logic_vector(22 downto 0); -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                               : std_logic;                     -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                         : std_logic;                     -- limiter:rsp_src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                               : std_logic;                     -- limiter:rsp_src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                       : std_logic;                     -- limiter:rsp_src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                                : std_logic_vector(97 downto 0); -- limiter:rsp_src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                             : std_logic_vector(22 downto 0); -- limiter:rsp_src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                               : std_logic;                     -- nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal addr_router_001_src_endofpacket                                                                     : std_logic;                     -- addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	signal addr_router_001_src_valid                                                                           : std_logic;                     -- addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	signal addr_router_001_src_startofpacket                                                                   : std_logic;                     -- addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	signal addr_router_001_src_data                                                                            : std_logic_vector(97 downto 0); -- addr_router_001:src_data -> limiter_001:cmd_sink_data
	signal addr_router_001_src_channel                                                                         : std_logic_vector(22 downto 0); -- addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	signal addr_router_001_src_ready                                                                           : std_logic;                     -- limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	signal limiter_001_rsp_src_endofpacket                                                                     : std_logic;                     -- limiter_001:rsp_src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_001_rsp_src_valid                                                                           : std_logic;                     -- limiter_001:rsp_src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_001_rsp_src_startofpacket                                                                   : std_logic;                     -- limiter_001:rsp_src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_001_rsp_src_data                                                                            : std_logic_vector(97 downto 0); -- limiter_001:rsp_src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_001_rsp_src_channel                                                                         : std_logic_vector(22 downto 0); -- limiter_001:rsp_src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_001_rsp_src_ready                                                                           : std_logic;                     -- nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                                   : std_logic;                     -- burst_adapter:source0_endofpacket -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                         : std_logic;                     -- burst_adapter:source0_valid -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                 : std_logic;                     -- burst_adapter:source0_startofpacket -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                          : std_logic_vector(79 downto 0); -- burst_adapter:source0_data -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                         : std_logic;                     -- SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                       : std_logic_vector(22 downto 0); -- burst_adapter:source0_channel -> SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                               : std_logic;                     -- burst_adapter_001:source0_endofpacket -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                     : std_logic;                     -- burst_adapter_001:source0_valid -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                             : std_logic;                     -- burst_adapter_001:source0_startofpacket -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                      : std_logic_vector(79 downto 0); -- burst_adapter_001:source0_data -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                     : std_logic;                     -- AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                   : std_logic_vector(22 downto 0); -- burst_adapter_001:source0_channel -> AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                      : std_logic;                     -- rst_controller:reset_out -> [AUDIO_DAC_FIFO_0_s0_translator:reset, AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent:reset, AUDIO_DAC_FIFO_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SRAM_DE2_0_s0_translator:reset, SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent:reset, SRAM_DE2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, audio_sos_s1_translator:reset, audio_sos_s1_translator_avalon_universal_slave_0_agent:reset, audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter:reset, burst_adapter_001:reset, clap_irq_s1_translator:reset, clap_irq_s1_translator_avalon_universal_slave_0_agent:reset, clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_011:reset, cmd_xbar_mux_012:reset, cmd_xbar_mux_013:reset, cmd_xbar_mux_014:reset, cmd_xbar_mux_015:reset, cmd_xbar_mux_016:reset, cmd_xbar_mux_017:reset, cmd_xbar_mux_018:reset, cmd_xbar_mux_019:reset, color_out_s1_translator:reset, color_out_s1_translator_avalon_universal_slave_0_agent:reset, color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dac_irq_s1_translator:reset, dac_irq_s1_translator_avalon_universal_slave_0_agent:reset, dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, hh_irq_s1_translator:reset, hh_irq_s1_translator_avalon_universal_slave_0_agent:reset, hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, in_bus_s1_translator:reset, in_bus_s1_translator_avalon_universal_slave_0_agent:reset, in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, irq_mapper:reset, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, kb_data_s1_translator:reset, kb_data_s1_translator_avalon_universal_slave_0_agent:reset, kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, kb_irq_s1_translator:reset, kb_irq_s1_translator_avalon_universal_slave_0_agent:reset, kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, kick_irq_s1_translator:reset, kick_irq_s1_translator_avalon_universal_slave_0_agent:reset, kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_r_s1_translator:reset, led_r_s1_translator_avalon_universal_slave_0_agent:reset, led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, seq_clap_s1_translator:reset, seq_clap_s1_translator_avalon_universal_slave_0_agent:reset, seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, seq_hh_s1_translator:reset, seq_hh_s1_translator_avalon_universal_slave_0_agent:reset, seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, seq_kick_s1_translator:reset, seq_kick_s1_translator_avalon_universal_slave_0_agent:reset, seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, seq_snare_s1_translator:reset, seq_snare_s1_translator_avalon_universal_slave_0_agent:reset, seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, snare_irq_s1_translator:reset, snare_irq_s1_translator_avalon_universal_slave_0_agent:reset, snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, wr_address_s1_translator:reset, wr_address_s1_translator_avalon_universal_slave_0_agent:reset, wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, wr_en_s1_translator:reset, wr_en_s1_translator_avalon_universal_slave_0_agent:reset, wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal nios2_qsys_0_jtag_debug_module_reset_reset                                                          : std_logic;                     -- nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	signal cmd_xbar_demux_src0_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                           : std_logic;                     -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                           : std_logic;                     -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                           : std_logic;                     -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_src3_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                           : std_logic;                     -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_src4_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal cmd_xbar_demux_src4_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	signal cmd_xbar_demux_src4_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	signal cmd_xbar_demux_src4_ready                                                                           : std_logic;                     -- cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	signal cmd_xbar_demux_src5_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	signal cmd_xbar_demux_src5_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	signal cmd_xbar_demux_src5_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	signal cmd_xbar_demux_src5_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	signal cmd_xbar_demux_src5_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	signal cmd_xbar_demux_src5_ready                                                                           : std_logic;                     -- cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	signal cmd_xbar_demux_src6_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src6_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	signal cmd_xbar_demux_src6_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src6_valid -> cmd_xbar_mux_006:sink0_valid
	signal cmd_xbar_demux_src6_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src6_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	signal cmd_xbar_demux_src6_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src6_data -> cmd_xbar_mux_006:sink0_data
	signal cmd_xbar_demux_src6_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src6_channel -> cmd_xbar_mux_006:sink0_channel
	signal cmd_xbar_demux_src6_ready                                                                           : std_logic;                     -- cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux:src6_ready
	signal cmd_xbar_demux_src7_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	signal cmd_xbar_demux_src7_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	signal cmd_xbar_demux_src7_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	signal cmd_xbar_demux_src7_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	signal cmd_xbar_demux_src7_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	signal cmd_xbar_demux_src7_ready                                                                           : std_logic;                     -- cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	signal cmd_xbar_demux_src8_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	signal cmd_xbar_demux_src8_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	signal cmd_xbar_demux_src8_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	signal cmd_xbar_demux_src8_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	signal cmd_xbar_demux_src8_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	signal cmd_xbar_demux_src8_ready                                                                           : std_logic;                     -- cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	signal cmd_xbar_demux_src9_endofpacket                                                                     : std_logic;                     -- cmd_xbar_demux:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	signal cmd_xbar_demux_src9_valid                                                                           : std_logic;                     -- cmd_xbar_demux:src9_valid -> cmd_xbar_mux_009:sink0_valid
	signal cmd_xbar_demux_src9_startofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	signal cmd_xbar_demux_src9_data                                                                            : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src9_data -> cmd_xbar_mux_009:sink0_data
	signal cmd_xbar_demux_src9_channel                                                                         : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src9_channel -> cmd_xbar_mux_009:sink0_channel
	signal cmd_xbar_demux_src9_ready                                                                           : std_logic;                     -- cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux:src9_ready
	signal cmd_xbar_demux_src10_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	signal cmd_xbar_demux_src10_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src10_valid -> cmd_xbar_mux_010:sink0_valid
	signal cmd_xbar_demux_src10_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	signal cmd_xbar_demux_src10_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src10_data -> cmd_xbar_mux_010:sink0_data
	signal cmd_xbar_demux_src10_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src10_channel -> cmd_xbar_mux_010:sink0_channel
	signal cmd_xbar_demux_src10_ready                                                                          : std_logic;                     -- cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux:src10_ready
	signal cmd_xbar_demux_src11_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src11_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	signal cmd_xbar_demux_src11_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src11_valid -> cmd_xbar_mux_011:sink0_valid
	signal cmd_xbar_demux_src11_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src11_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	signal cmd_xbar_demux_src11_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src11_data -> cmd_xbar_mux_011:sink0_data
	signal cmd_xbar_demux_src11_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src11_channel -> cmd_xbar_mux_011:sink0_channel
	signal cmd_xbar_demux_src11_ready                                                                          : std_logic;                     -- cmd_xbar_mux_011:sink0_ready -> cmd_xbar_demux:src11_ready
	signal cmd_xbar_demux_src12_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src12_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	signal cmd_xbar_demux_src12_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src12_valid -> cmd_xbar_mux_012:sink0_valid
	signal cmd_xbar_demux_src12_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src12_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	signal cmd_xbar_demux_src12_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src12_data -> cmd_xbar_mux_012:sink0_data
	signal cmd_xbar_demux_src12_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src12_channel -> cmd_xbar_mux_012:sink0_channel
	signal cmd_xbar_demux_src12_ready                                                                          : std_logic;                     -- cmd_xbar_mux_012:sink0_ready -> cmd_xbar_demux:src12_ready
	signal cmd_xbar_demux_src13_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	signal cmd_xbar_demux_src13_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src13_valid -> cmd_xbar_mux_013:sink0_valid
	signal cmd_xbar_demux_src13_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	signal cmd_xbar_demux_src13_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src13_data -> cmd_xbar_mux_013:sink0_data
	signal cmd_xbar_demux_src13_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src13_channel -> cmd_xbar_mux_013:sink0_channel
	signal cmd_xbar_demux_src13_ready                                                                          : std_logic;                     -- cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux:src13_ready
	signal cmd_xbar_demux_src14_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src14_endofpacket -> cmd_xbar_mux_014:sink0_endofpacket
	signal cmd_xbar_demux_src14_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src14_valid -> cmd_xbar_mux_014:sink0_valid
	signal cmd_xbar_demux_src14_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src14_startofpacket -> cmd_xbar_mux_014:sink0_startofpacket
	signal cmd_xbar_demux_src14_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src14_data -> cmd_xbar_mux_014:sink0_data
	signal cmd_xbar_demux_src14_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src14_channel -> cmd_xbar_mux_014:sink0_channel
	signal cmd_xbar_demux_src14_ready                                                                          : std_logic;                     -- cmd_xbar_mux_014:sink0_ready -> cmd_xbar_demux:src14_ready
	signal cmd_xbar_demux_src15_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src15_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	signal cmd_xbar_demux_src15_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src15_valid -> cmd_xbar_mux_015:sink0_valid
	signal cmd_xbar_demux_src15_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src15_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	signal cmd_xbar_demux_src15_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src15_data -> cmd_xbar_mux_015:sink0_data
	signal cmd_xbar_demux_src15_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src15_channel -> cmd_xbar_mux_015:sink0_channel
	signal cmd_xbar_demux_src15_ready                                                                          : std_logic;                     -- cmd_xbar_mux_015:sink0_ready -> cmd_xbar_demux:src15_ready
	signal cmd_xbar_demux_src16_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src16_endofpacket -> cmd_xbar_mux_016:sink0_endofpacket
	signal cmd_xbar_demux_src16_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src16_valid -> cmd_xbar_mux_016:sink0_valid
	signal cmd_xbar_demux_src16_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src16_startofpacket -> cmd_xbar_mux_016:sink0_startofpacket
	signal cmd_xbar_demux_src16_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src16_data -> cmd_xbar_mux_016:sink0_data
	signal cmd_xbar_demux_src16_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src16_channel -> cmd_xbar_mux_016:sink0_channel
	signal cmd_xbar_demux_src16_ready                                                                          : std_logic;                     -- cmd_xbar_mux_016:sink0_ready -> cmd_xbar_demux:src16_ready
	signal cmd_xbar_demux_src17_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src17_endofpacket -> cmd_xbar_mux_017:sink0_endofpacket
	signal cmd_xbar_demux_src17_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src17_valid -> cmd_xbar_mux_017:sink0_valid
	signal cmd_xbar_demux_src17_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src17_startofpacket -> cmd_xbar_mux_017:sink0_startofpacket
	signal cmd_xbar_demux_src17_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src17_data -> cmd_xbar_mux_017:sink0_data
	signal cmd_xbar_demux_src17_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src17_channel -> cmd_xbar_mux_017:sink0_channel
	signal cmd_xbar_demux_src17_ready                                                                          : std_logic;                     -- cmd_xbar_mux_017:sink0_ready -> cmd_xbar_demux:src17_ready
	signal cmd_xbar_demux_src18_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src18_endofpacket -> cmd_xbar_mux_018:sink0_endofpacket
	signal cmd_xbar_demux_src18_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src18_valid -> cmd_xbar_mux_018:sink0_valid
	signal cmd_xbar_demux_src18_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src18_startofpacket -> cmd_xbar_mux_018:sink0_startofpacket
	signal cmd_xbar_demux_src18_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src18_data -> cmd_xbar_mux_018:sink0_data
	signal cmd_xbar_demux_src18_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src18_channel -> cmd_xbar_mux_018:sink0_channel
	signal cmd_xbar_demux_src18_ready                                                                          : std_logic;                     -- cmd_xbar_mux_018:sink0_ready -> cmd_xbar_demux:src18_ready
	signal cmd_xbar_demux_src19_endofpacket                                                                    : std_logic;                     -- cmd_xbar_demux:src19_endofpacket -> cmd_xbar_mux_019:sink0_endofpacket
	signal cmd_xbar_demux_src19_valid                                                                          : std_logic;                     -- cmd_xbar_demux:src19_valid -> cmd_xbar_mux_019:sink0_valid
	signal cmd_xbar_demux_src19_startofpacket                                                                  : std_logic;                     -- cmd_xbar_demux:src19_startofpacket -> cmd_xbar_mux_019:sink0_startofpacket
	signal cmd_xbar_demux_src19_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_demux:src19_data -> cmd_xbar_mux_019:sink0_data
	signal cmd_xbar_demux_src19_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_demux:src19_channel -> cmd_xbar_mux_019:sink0_channel
	signal cmd_xbar_demux_src19_ready                                                                          : std_logic;                     -- cmd_xbar_mux_019:sink0_ready -> cmd_xbar_demux:src19_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                       : std_logic;                     -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                       : std_logic;                     -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                       : std_logic;                     -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src3_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src3_ready                                                                       : std_logic;                     -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	signal cmd_xbar_demux_001_src4_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	signal cmd_xbar_demux_001_src4_ready                                                                       : std_logic;                     -- cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	signal cmd_xbar_demux_001_src5_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	signal cmd_xbar_demux_001_src5_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	signal cmd_xbar_demux_001_src5_ready                                                                       : std_logic;                     -- cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	signal cmd_xbar_demux_001_src6_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src6_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src6_valid -> cmd_xbar_mux_006:sink1_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src6_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src6_data -> cmd_xbar_mux_006:sink1_data
	signal cmd_xbar_demux_001_src6_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src6_channel -> cmd_xbar_mux_006:sink1_channel
	signal cmd_xbar_demux_001_src6_ready                                                                       : std_logic;                     -- cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_001:src6_ready
	signal cmd_xbar_demux_001_src7_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	signal cmd_xbar_demux_001_src7_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	signal cmd_xbar_demux_001_src7_ready                                                                       : std_logic;                     -- cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	signal cmd_xbar_demux_001_src8_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink1_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink1_data
	signal cmd_xbar_demux_001_src8_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink1_channel
	signal cmd_xbar_demux_001_src8_ready                                                                       : std_logic;                     -- cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src8_ready
	signal cmd_xbar_demux_001_src9_endofpacket                                                                 : std_logic;                     -- cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                       : std_logic;                     -- cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink1_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                        : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink1_data
	signal cmd_xbar_demux_001_src9_channel                                                                     : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink1_channel
	signal cmd_xbar_demux_001_src9_ready                                                                       : std_logic;                     -- cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_001:src9_ready
	signal cmd_xbar_demux_001_src10_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink1_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink1_data
	signal cmd_xbar_demux_001_src10_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink1_channel
	signal cmd_xbar_demux_001_src10_ready                                                                      : std_logic;                     -- cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_001:src10_ready
	signal cmd_xbar_demux_001_src11_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src11_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	signal cmd_xbar_demux_001_src11_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src11_valid -> cmd_xbar_mux_011:sink1_valid
	signal cmd_xbar_demux_001_src11_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src11_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	signal cmd_xbar_demux_001_src11_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src11_data -> cmd_xbar_mux_011:sink1_data
	signal cmd_xbar_demux_001_src11_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src11_channel -> cmd_xbar_mux_011:sink1_channel
	signal cmd_xbar_demux_001_src11_ready                                                                      : std_logic;                     -- cmd_xbar_mux_011:sink1_ready -> cmd_xbar_demux_001:src11_ready
	signal cmd_xbar_demux_001_src12_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src12_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	signal cmd_xbar_demux_001_src12_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src12_valid -> cmd_xbar_mux_012:sink1_valid
	signal cmd_xbar_demux_001_src12_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src12_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	signal cmd_xbar_demux_001_src12_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src12_data -> cmd_xbar_mux_012:sink1_data
	signal cmd_xbar_demux_001_src12_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src12_channel -> cmd_xbar_mux_012:sink1_channel
	signal cmd_xbar_demux_001_src12_ready                                                                      : std_logic;                     -- cmd_xbar_mux_012:sink1_ready -> cmd_xbar_demux_001:src12_ready
	signal cmd_xbar_demux_001_src13_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src13_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	signal cmd_xbar_demux_001_src13_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src13_valid -> cmd_xbar_mux_013:sink1_valid
	signal cmd_xbar_demux_001_src13_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src13_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	signal cmd_xbar_demux_001_src13_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src13_data -> cmd_xbar_mux_013:sink1_data
	signal cmd_xbar_demux_001_src13_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src13_channel -> cmd_xbar_mux_013:sink1_channel
	signal cmd_xbar_demux_001_src13_ready                                                                      : std_logic;                     -- cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_001:src13_ready
	signal cmd_xbar_demux_001_src14_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src14_endofpacket -> cmd_xbar_mux_014:sink1_endofpacket
	signal cmd_xbar_demux_001_src14_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src14_valid -> cmd_xbar_mux_014:sink1_valid
	signal cmd_xbar_demux_001_src14_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src14_startofpacket -> cmd_xbar_mux_014:sink1_startofpacket
	signal cmd_xbar_demux_001_src14_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src14_data -> cmd_xbar_mux_014:sink1_data
	signal cmd_xbar_demux_001_src14_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src14_channel -> cmd_xbar_mux_014:sink1_channel
	signal cmd_xbar_demux_001_src14_ready                                                                      : std_logic;                     -- cmd_xbar_mux_014:sink1_ready -> cmd_xbar_demux_001:src14_ready
	signal cmd_xbar_demux_001_src15_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src15_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	signal cmd_xbar_demux_001_src15_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src15_valid -> cmd_xbar_mux_015:sink1_valid
	signal cmd_xbar_demux_001_src15_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src15_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	signal cmd_xbar_demux_001_src15_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src15_data -> cmd_xbar_mux_015:sink1_data
	signal cmd_xbar_demux_001_src15_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src15_channel -> cmd_xbar_mux_015:sink1_channel
	signal cmd_xbar_demux_001_src15_ready                                                                      : std_logic;                     -- cmd_xbar_mux_015:sink1_ready -> cmd_xbar_demux_001:src15_ready
	signal cmd_xbar_demux_001_src16_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src16_endofpacket -> cmd_xbar_mux_016:sink1_endofpacket
	signal cmd_xbar_demux_001_src16_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src16_valid -> cmd_xbar_mux_016:sink1_valid
	signal cmd_xbar_demux_001_src16_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src16_startofpacket -> cmd_xbar_mux_016:sink1_startofpacket
	signal cmd_xbar_demux_001_src16_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src16_data -> cmd_xbar_mux_016:sink1_data
	signal cmd_xbar_demux_001_src16_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src16_channel -> cmd_xbar_mux_016:sink1_channel
	signal cmd_xbar_demux_001_src16_ready                                                                      : std_logic;                     -- cmd_xbar_mux_016:sink1_ready -> cmd_xbar_demux_001:src16_ready
	signal cmd_xbar_demux_001_src17_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src17_endofpacket -> cmd_xbar_mux_017:sink1_endofpacket
	signal cmd_xbar_demux_001_src17_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src17_valid -> cmd_xbar_mux_017:sink1_valid
	signal cmd_xbar_demux_001_src17_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src17_startofpacket -> cmd_xbar_mux_017:sink1_startofpacket
	signal cmd_xbar_demux_001_src17_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src17_data -> cmd_xbar_mux_017:sink1_data
	signal cmd_xbar_demux_001_src17_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src17_channel -> cmd_xbar_mux_017:sink1_channel
	signal cmd_xbar_demux_001_src17_ready                                                                      : std_logic;                     -- cmd_xbar_mux_017:sink1_ready -> cmd_xbar_demux_001:src17_ready
	signal cmd_xbar_demux_001_src18_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src18_endofpacket -> cmd_xbar_mux_018:sink1_endofpacket
	signal cmd_xbar_demux_001_src18_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src18_valid -> cmd_xbar_mux_018:sink1_valid
	signal cmd_xbar_demux_001_src18_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src18_startofpacket -> cmd_xbar_mux_018:sink1_startofpacket
	signal cmd_xbar_demux_001_src18_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src18_data -> cmd_xbar_mux_018:sink1_data
	signal cmd_xbar_demux_001_src18_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src18_channel -> cmd_xbar_mux_018:sink1_channel
	signal cmd_xbar_demux_001_src18_ready                                                                      : std_logic;                     -- cmd_xbar_mux_018:sink1_ready -> cmd_xbar_demux_001:src18_ready
	signal cmd_xbar_demux_001_src19_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src19_endofpacket -> cmd_xbar_mux_019:sink1_endofpacket
	signal cmd_xbar_demux_001_src19_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src19_valid -> cmd_xbar_mux_019:sink1_valid
	signal cmd_xbar_demux_001_src19_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src19_startofpacket -> cmd_xbar_mux_019:sink1_startofpacket
	signal cmd_xbar_demux_001_src19_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src19_data -> cmd_xbar_mux_019:sink1_data
	signal cmd_xbar_demux_001_src19_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src19_channel -> cmd_xbar_mux_019:sink1_channel
	signal cmd_xbar_demux_001_src19_ready                                                                      : std_logic;                     -- cmd_xbar_mux_019:sink1_ready -> cmd_xbar_demux_001:src19_ready
	signal cmd_xbar_demux_001_src20_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src20_endofpacket -> kb_data_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src20_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src20_valid -> kb_data_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src20_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src20_startofpacket -> kb_data_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src20_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src20_data -> kb_data_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src20_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src20_channel -> kb_data_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src21_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src21_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_demux_001_src21_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src21_valid -> width_adapter_002:in_valid
	signal cmd_xbar_demux_001_src21_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src21_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_demux_001_src21_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src21_data -> width_adapter_002:in_data
	signal cmd_xbar_demux_001_src21_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src21_channel -> width_adapter_002:in_channel
	signal cmd_xbar_demux_001_src22_endofpacket                                                                : std_logic;                     -- cmd_xbar_demux_001:src22_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src22_valid                                                                      : std_logic;                     -- cmd_xbar_demux_001:src22_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src22_startofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src22_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src22_data                                                                       : std_logic_vector(97 downto 0); -- cmd_xbar_demux_001:src22_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src22_channel                                                                    : std_logic_vector(22 downto 0); -- cmd_xbar_demux_001:src22_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                     : std_logic;                     -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                           : std_logic;                     -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                   : std_logic;                     -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                            : std_logic_vector(97 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                         : std_logic_vector(22 downto 0); -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                           : std_logic;                     -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                     : std_logic;                     -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                           : std_logic;                     -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                   : std_logic;                     -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                            : std_logic_vector(97 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                         : std_logic_vector(22 downto 0); -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                           : std_logic;                     -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_004_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_005_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_006_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src1_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_007_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_008_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src1_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_009_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src1_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_010_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal rsp_xbar_demux_010_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_001:sink10_valid
	signal rsp_xbar_demux_010_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal rsp_xbar_demux_010_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_001:sink10_data
	signal rsp_xbar_demux_010_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_001:sink10_channel
	signal rsp_xbar_demux_010_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src1_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_011_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_011:src1_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	signal rsp_xbar_demux_011_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_011:src1_valid -> rsp_xbar_mux_001:sink11_valid
	signal rsp_xbar_demux_011_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_011:src1_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	signal rsp_xbar_demux_011_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_011:src1_data -> rsp_xbar_mux_001:sink11_data
	signal rsp_xbar_demux_011_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_011:src1_channel -> rsp_xbar_mux_001:sink11_channel
	signal rsp_xbar_demux_011_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src1_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_012_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_012:src1_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	signal rsp_xbar_demux_012_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_012:src1_valid -> rsp_xbar_mux_001:sink12_valid
	signal rsp_xbar_demux_012_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_012:src1_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	signal rsp_xbar_demux_012_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_012:src1_data -> rsp_xbar_mux_001:sink12_data
	signal rsp_xbar_demux_012_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_012:src1_channel -> rsp_xbar_mux_001:sink12_channel
	signal rsp_xbar_demux_012_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src1_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_013_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	signal rsp_xbar_demux_013_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_001:sink13_valid
	signal rsp_xbar_demux_013_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	signal rsp_xbar_demux_013_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_001:sink13_data
	signal rsp_xbar_demux_013_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_001:sink13_channel
	signal rsp_xbar_demux_013_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src1_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	signal rsp_xbar_demux_014_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	signal rsp_xbar_demux_014_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	signal rsp_xbar_demux_014_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_014:src1_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	signal rsp_xbar_demux_014_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_014:src1_valid -> rsp_xbar_mux_001:sink14_valid
	signal rsp_xbar_demux_014_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_014:src1_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	signal rsp_xbar_demux_014_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_014:src1_data -> rsp_xbar_mux_001:sink14_data
	signal rsp_xbar_demux_014_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_014:src1_channel -> rsp_xbar_mux_001:sink14_channel
	signal rsp_xbar_demux_014_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src1_ready
	signal rsp_xbar_demux_015_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	signal rsp_xbar_demux_015_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux:sink15_valid
	signal rsp_xbar_demux_015_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	signal rsp_xbar_demux_015_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_015:src0_data -> rsp_xbar_mux:sink15_data
	signal rsp_xbar_demux_015_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux:sink15_channel
	signal rsp_xbar_demux_015_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink15_ready -> rsp_xbar_demux_015:src0_ready
	signal rsp_xbar_demux_015_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_015:src1_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	signal rsp_xbar_demux_015_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_015:src1_valid -> rsp_xbar_mux_001:sink15_valid
	signal rsp_xbar_demux_015_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_015:src1_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	signal rsp_xbar_demux_015_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_015:src1_data -> rsp_xbar_mux_001:sink15_data
	signal rsp_xbar_demux_015_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_015:src1_channel -> rsp_xbar_mux_001:sink15_channel
	signal rsp_xbar_demux_015_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src1_ready
	signal rsp_xbar_demux_016_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux:sink16_endofpacket
	signal rsp_xbar_demux_016_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux:sink16_valid
	signal rsp_xbar_demux_016_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux:sink16_startofpacket
	signal rsp_xbar_demux_016_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_016:src0_data -> rsp_xbar_mux:sink16_data
	signal rsp_xbar_demux_016_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux:sink16_channel
	signal rsp_xbar_demux_016_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink16_ready -> rsp_xbar_demux_016:src0_ready
	signal rsp_xbar_demux_016_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_016:src1_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	signal rsp_xbar_demux_016_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_016:src1_valid -> rsp_xbar_mux_001:sink16_valid
	signal rsp_xbar_demux_016_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_016:src1_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	signal rsp_xbar_demux_016_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_016:src1_data -> rsp_xbar_mux_001:sink16_data
	signal rsp_xbar_demux_016_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_016:src1_channel -> rsp_xbar_mux_001:sink16_channel
	signal rsp_xbar_demux_016_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src1_ready
	signal rsp_xbar_demux_017_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux:sink17_endofpacket
	signal rsp_xbar_demux_017_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux:sink17_valid
	signal rsp_xbar_demux_017_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux:sink17_startofpacket
	signal rsp_xbar_demux_017_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_017:src0_data -> rsp_xbar_mux:sink17_data
	signal rsp_xbar_demux_017_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux:sink17_channel
	signal rsp_xbar_demux_017_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink17_ready -> rsp_xbar_demux_017:src0_ready
	signal rsp_xbar_demux_017_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_017:src1_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	signal rsp_xbar_demux_017_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_017:src1_valid -> rsp_xbar_mux_001:sink17_valid
	signal rsp_xbar_demux_017_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_017:src1_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	signal rsp_xbar_demux_017_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_017:src1_data -> rsp_xbar_mux_001:sink17_data
	signal rsp_xbar_demux_017_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_017:src1_channel -> rsp_xbar_mux_001:sink17_channel
	signal rsp_xbar_demux_017_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src1_ready
	signal rsp_xbar_demux_018_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux:sink18_endofpacket
	signal rsp_xbar_demux_018_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux:sink18_valid
	signal rsp_xbar_demux_018_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux:sink18_startofpacket
	signal rsp_xbar_demux_018_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_018:src0_data -> rsp_xbar_mux:sink18_data
	signal rsp_xbar_demux_018_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux:sink18_channel
	signal rsp_xbar_demux_018_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink18_ready -> rsp_xbar_demux_018:src0_ready
	signal rsp_xbar_demux_018_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_018:src1_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	signal rsp_xbar_demux_018_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_018:src1_valid -> rsp_xbar_mux_001:sink18_valid
	signal rsp_xbar_demux_018_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_018:src1_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	signal rsp_xbar_demux_018_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_018:src1_data -> rsp_xbar_mux_001:sink18_data
	signal rsp_xbar_demux_018_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_018:src1_channel -> rsp_xbar_mux_001:sink18_channel
	signal rsp_xbar_demux_018_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src1_ready
	signal rsp_xbar_demux_019_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux:sink19_endofpacket
	signal rsp_xbar_demux_019_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux:sink19_valid
	signal rsp_xbar_demux_019_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux:sink19_startofpacket
	signal rsp_xbar_demux_019_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_019:src0_data -> rsp_xbar_mux:sink19_data
	signal rsp_xbar_demux_019_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux:sink19_channel
	signal rsp_xbar_demux_019_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux:sink19_ready -> rsp_xbar_demux_019:src0_ready
	signal rsp_xbar_demux_019_src1_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_019:src1_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	signal rsp_xbar_demux_019_src1_valid                                                                       : std_logic;                     -- rsp_xbar_demux_019:src1_valid -> rsp_xbar_mux_001:sink19_valid
	signal rsp_xbar_demux_019_src1_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_019:src1_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	signal rsp_xbar_demux_019_src1_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_019:src1_data -> rsp_xbar_mux_001:sink19_data
	signal rsp_xbar_demux_019_src1_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_019:src1_channel -> rsp_xbar_mux_001:sink19_channel
	signal rsp_xbar_demux_019_src1_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src1_ready
	signal rsp_xbar_demux_020_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	signal rsp_xbar_demux_020_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	signal rsp_xbar_demux_020_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	signal rsp_xbar_demux_020_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	signal rsp_xbar_demux_020_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	signal rsp_xbar_demux_020_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	signal rsp_xbar_demux_021_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	signal rsp_xbar_demux_021_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	signal rsp_xbar_demux_021_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	signal rsp_xbar_demux_021_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	signal rsp_xbar_demux_021_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	signal rsp_xbar_demux_021_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	signal rsp_xbar_demux_022_src0_endofpacket                                                                 : std_logic;                     -- rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	signal rsp_xbar_demux_022_src0_valid                                                                       : std_logic;                     -- rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	signal rsp_xbar_demux_022_src0_startofpacket                                                               : std_logic;                     -- rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	signal rsp_xbar_demux_022_src0_data                                                                        : std_logic_vector(97 downto 0); -- rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	signal rsp_xbar_demux_022_src0_channel                                                                     : std_logic_vector(22 downto 0); -- rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	signal rsp_xbar_demux_022_src0_ready                                                                       : std_logic;                     -- rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	signal limiter_cmd_src_endofpacket                                                                         : std_logic;                     -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                       : std_logic;                     -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                                : std_logic_vector(97 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                             : std_logic_vector(22 downto 0); -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                               : std_logic;                     -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                        : std_logic;                     -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                              : std_logic;                     -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                                      : std_logic;                     -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                               : std_logic_vector(97 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                            : std_logic_vector(22 downto 0); -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                              : std_logic;                     -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal limiter_001_cmd_src_endofpacket                                                                     : std_logic;                     -- limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal limiter_001_cmd_src_startofpacket                                                                   : std_logic;                     -- limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal limiter_001_cmd_src_data                                                                            : std_logic_vector(97 downto 0); -- limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	signal limiter_001_cmd_src_channel                                                                         : std_logic_vector(22 downto 0); -- limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	signal limiter_001_cmd_src_ready                                                                           : std_logic;                     -- cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                    : std_logic;                     -- rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                          : std_logic;                     -- rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                  : std_logic;                     -- rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                           : std_logic_vector(97 downto 0); -- rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	signal rsp_xbar_mux_001_src_channel                                                                        : std_logic_vector(22 downto 0); -- rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	signal rsp_xbar_mux_001_src_ready                                                                          : std_logic;                     -- limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                        : std_logic;                     -- cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                              : std_logic;                     -- cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                      : std_logic;                     -- cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                               : std_logic_vector(97 downto 0); -- cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                            : std_logic_vector(22 downto 0); -- cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                              : std_logic;                     -- nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                           : std_logic;                     -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                 : std_logic;                     -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                         : std_logic;                     -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                  : std_logic_vector(97 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                               : std_logic_vector(22 downto 0); -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                 : std_logic;                     -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_002:src_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_002:src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_002:src_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_002:src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_002_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_002:src_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_002_src_ready                                                                          : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                                       : std_logic;                     -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                             : std_logic;                     -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                     : std_logic;                     -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_mux_003_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_003:src_endofpacket -> audio_sos_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_003:src_valid -> audio_sos_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_003:src_startofpacket -> audio_sos_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_003:src_data -> audio_sos_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_003_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_003:src_channel -> audio_sos_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_003_src_ready                                                                          : std_logic;                     -- audio_sos_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	signal id_router_003_src_endofpacket                                                                       : std_logic;                     -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                             : std_logic;                     -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                     : std_logic;                     -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_004:src_endofpacket -> dac_irq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_004:src_valid -> dac_irq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_004:src_startofpacket -> dac_irq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_004:src_data -> dac_irq_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_004_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_004:src_channel -> dac_irq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_004_src_ready                                                                          : std_logic;                     -- dac_irq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                       : std_logic;                     -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                             : std_logic;                     -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                     : std_logic;                     -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_mux_005_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_005:src_endofpacket -> clap_irq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_005_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_005:src_valid -> clap_irq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_005_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_005:src_startofpacket -> clap_irq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_005_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_005:src_data -> clap_irq_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_005_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_005:src_channel -> clap_irq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_005_src_ready                                                                          : std_logic;                     -- clap_irq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	signal id_router_005_src_endofpacket                                                                       : std_logic;                     -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                             : std_logic;                     -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                     : std_logic;                     -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_mux_006_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_006:src_endofpacket -> hh_irq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_006_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_006:src_valid -> hh_irq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_006_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_006:src_startofpacket -> hh_irq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_006_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_006:src_data -> hh_irq_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_006_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_006:src_channel -> hh_irq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_006_src_ready                                                                          : std_logic;                     -- hh_irq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_006:src_ready
	signal id_router_006_src_endofpacket                                                                       : std_logic;                     -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                             : std_logic;                     -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                     : std_logic;                     -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_mux_007_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_007:src_endofpacket -> snare_irq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_007_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_007:src_valid -> snare_irq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_007_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_007:src_startofpacket -> snare_irq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_007_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_007:src_data -> snare_irq_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_007_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_007:src_channel -> snare_irq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_007_src_ready                                                                          : std_logic;                     -- snare_irq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	signal id_router_007_src_endofpacket                                                                       : std_logic;                     -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                             : std_logic;                     -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                     : std_logic;                     -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_mux_008_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_008:src_endofpacket -> kick_irq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_008_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_008:src_valid -> kick_irq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_008_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_008:src_startofpacket -> kick_irq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_008_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_008:src_data -> kick_irq_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_008_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_008:src_channel -> kick_irq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_008_src_ready                                                                          : std_logic;                     -- kick_irq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	signal id_router_008_src_endofpacket                                                                       : std_logic;                     -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                             : std_logic;                     -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                     : std_logic;                     -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_mux_009_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_009:src_endofpacket -> kb_irq_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_009_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_009:src_valid -> kb_irq_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_009_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_009:src_startofpacket -> kb_irq_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_009_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_009:src_data -> kb_irq_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_009_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_009:src_channel -> kb_irq_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_009_src_ready                                                                          : std_logic;                     -- kb_irq_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	signal id_router_009_src_endofpacket                                                                       : std_logic;                     -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                             : std_logic;                     -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                     : std_logic;                     -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_mux_010_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_010:src_endofpacket -> seq_hh_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_010_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_010:src_valid -> seq_hh_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_010_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_010:src_startofpacket -> seq_hh_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_010_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_010:src_data -> seq_hh_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_010_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_010:src_channel -> seq_hh_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_010_src_ready                                                                          : std_logic;                     -- seq_hh_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	signal id_router_010_src_endofpacket                                                                       : std_logic;                     -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                             : std_logic;                     -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                     : std_logic;                     -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_mux_011_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_011:src_endofpacket -> seq_snare_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_011_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_011:src_valid -> seq_snare_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_011_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_011:src_startofpacket -> seq_snare_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_011_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_011:src_data -> seq_snare_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_011_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_011:src_channel -> seq_snare_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_011_src_ready                                                                          : std_logic;                     -- seq_snare_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_011:src_ready
	signal id_router_011_src_endofpacket                                                                       : std_logic;                     -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                             : std_logic;                     -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                     : std_logic;                     -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_mux_012_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_012:src_endofpacket -> led_r_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_012_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_012:src_valid -> led_r_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_012_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_012:src_startofpacket -> led_r_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_012_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_012:src_data -> led_r_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_012_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_012:src_channel -> led_r_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_012_src_ready                                                                          : std_logic;                     -- led_r_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_012:src_ready
	signal id_router_012_src_endofpacket                                                                       : std_logic;                     -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                             : std_logic;                     -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                     : std_logic;                     -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_mux_013_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_013:src_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_013_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_013:src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_013_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_013:src_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_013_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_013:src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_013_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_013:src_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_013_src_ready                                                                          : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	signal id_router_013_src_endofpacket                                                                       : std_logic;                     -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                             : std_logic;                     -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                                     : std_logic;                     -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal cmd_xbar_mux_014_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_014:src_endofpacket -> seq_clap_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_014_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_014:src_valid -> seq_clap_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_014_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_014:src_startofpacket -> seq_clap_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_014_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_014:src_data -> seq_clap_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_014_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_014:src_channel -> seq_clap_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_014_src_ready                                                                          : std_logic;                     -- seq_clap_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_014:src_ready
	signal id_router_014_src_endofpacket                                                                       : std_logic;                     -- id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal id_router_014_src_valid                                                                             : std_logic;                     -- id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	signal id_router_014_src_startofpacket                                                                     : std_logic;                     -- id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal id_router_014_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	signal id_router_014_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	signal id_router_014_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	signal cmd_xbar_mux_015_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_015:src_endofpacket -> seq_kick_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_015_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_015:src_valid -> seq_kick_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_015_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_015:src_startofpacket -> seq_kick_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_015_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_015:src_data -> seq_kick_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_015_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_015:src_channel -> seq_kick_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_015_src_ready                                                                          : std_logic;                     -- seq_kick_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_015:src_ready
	signal id_router_015_src_endofpacket                                                                       : std_logic;                     -- id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	signal id_router_015_src_valid                                                                             : std_logic;                     -- id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	signal id_router_015_src_startofpacket                                                                     : std_logic;                     -- id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	signal id_router_015_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	signal id_router_015_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	signal id_router_015_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	signal cmd_xbar_mux_016_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_016:src_endofpacket -> wr_address_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_016_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_016:src_valid -> wr_address_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_016_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_016:src_startofpacket -> wr_address_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_016_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_016:src_data -> wr_address_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_016_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_016:src_channel -> wr_address_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_016_src_ready                                                                          : std_logic;                     -- wr_address_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_016:src_ready
	signal id_router_016_src_endofpacket                                                                       : std_logic;                     -- id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	signal id_router_016_src_valid                                                                             : std_logic;                     -- id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	signal id_router_016_src_startofpacket                                                                     : std_logic;                     -- id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	signal id_router_016_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	signal id_router_016_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	signal id_router_016_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	signal cmd_xbar_mux_017_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_017:src_endofpacket -> color_out_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_017_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_017:src_valid -> color_out_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_017_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_017:src_startofpacket -> color_out_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_017_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_017:src_data -> color_out_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_017_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_017:src_channel -> color_out_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_017_src_ready                                                                          : std_logic;                     -- color_out_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_017:src_ready
	signal id_router_017_src_endofpacket                                                                       : std_logic;                     -- id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	signal id_router_017_src_valid                                                                             : std_logic;                     -- id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	signal id_router_017_src_startofpacket                                                                     : std_logic;                     -- id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	signal id_router_017_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	signal id_router_017_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	signal id_router_017_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	signal cmd_xbar_mux_018_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_018:src_endofpacket -> in_bus_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_018_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_018:src_valid -> in_bus_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_018_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_018:src_startofpacket -> in_bus_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_018_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_018:src_data -> in_bus_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_018_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_018:src_channel -> in_bus_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_018_src_ready                                                                          : std_logic;                     -- in_bus_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_018:src_ready
	signal id_router_018_src_endofpacket                                                                       : std_logic;                     -- id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	signal id_router_018_src_valid                                                                             : std_logic;                     -- id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	signal id_router_018_src_startofpacket                                                                     : std_logic;                     -- id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	signal id_router_018_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	signal id_router_018_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	signal id_router_018_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	signal cmd_xbar_mux_019_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_019:src_endofpacket -> wr_en_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_019_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_019:src_valid -> wr_en_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_019_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_019:src_startofpacket -> wr_en_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_019_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_019:src_data -> wr_en_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_019_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_019:src_channel -> wr_en_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_019_src_ready                                                                          : std_logic;                     -- wr_en_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_019:src_ready
	signal id_router_019_src_endofpacket                                                                       : std_logic;                     -- id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	signal id_router_019_src_valid                                                                             : std_logic;                     -- id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	signal id_router_019_src_startofpacket                                                                     : std_logic;                     -- id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	signal id_router_019_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	signal id_router_019_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	signal id_router_019_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	signal cmd_xbar_demux_001_src20_ready                                                                      : std_logic;                     -- kb_data_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	signal id_router_020_src_endofpacket                                                                       : std_logic;                     -- id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	signal id_router_020_src_valid                                                                             : std_logic;                     -- id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	signal id_router_020_src_startofpacket                                                                     : std_logic;                     -- id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	signal id_router_020_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	signal id_router_020_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	signal id_router_020_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	signal cmd_xbar_demux_001_src22_ready                                                                      : std_logic;                     -- timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	signal id_router_022_src_endofpacket                                                                       : std_logic;                     -- id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	signal id_router_022_src_valid                                                                             : std_logic;                     -- id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	signal id_router_022_src_startofpacket                                                                     : std_logic;                     -- id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	signal id_router_022_src_data                                                                              : std_logic_vector(97 downto 0); -- id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	signal id_router_022_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	signal id_router_022_src_ready                                                                             : std_logic;                     -- rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                    : std_logic;                     -- cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                          : std_logic;                     -- cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                           : std_logic_vector(97 downto 0); -- cmd_xbar_mux_001:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_001_src_channel                                                                        : std_logic_vector(22 downto 0); -- cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_001_src_ready                                                                          : std_logic;                     -- width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	signal width_adapter_src_endofpacket                                                                       : std_logic;                     -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                             : std_logic;                     -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                     : std_logic;                     -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                              : std_logic_vector(79 downto 0); -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                             : std_logic;                     -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                           : std_logic_vector(22 downto 0); -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_001_src_endofpacket                                                                       : std_logic;                     -- id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_001_src_valid                                                                             : std_logic;                     -- id_router_001:src_valid -> width_adapter_001:in_valid
	signal id_router_001_src_startofpacket                                                                     : std_logic;                     -- id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_001_src_data                                                                              : std_logic_vector(79 downto 0); -- id_router_001:src_data -> width_adapter_001:in_data
	signal id_router_001_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_001:src_channel -> width_adapter_001:in_channel
	signal id_router_001_src_ready                                                                             : std_logic;                     -- width_adapter_001:in_ready -> id_router_001:src_ready
	signal width_adapter_001_src_endofpacket                                                                   : std_logic;                     -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal width_adapter_001_src_valid                                                                         : std_logic;                     -- width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	signal width_adapter_001_src_startofpacket                                                                 : std_logic;                     -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal width_adapter_001_src_data                                                                          : std_logic_vector(97 downto 0); -- width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	signal width_adapter_001_src_ready                                                                         : std_logic;                     -- rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                       : std_logic_vector(22 downto 0); -- width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	signal cmd_xbar_demux_001_src21_ready                                                                      : std_logic;                     -- width_adapter_002:in_ready -> cmd_xbar_demux_001:src21_ready
	signal width_adapter_002_src_endofpacket                                                                   : std_logic;                     -- width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal width_adapter_002_src_valid                                                                         : std_logic;                     -- width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	signal width_adapter_002_src_startofpacket                                                                 : std_logic;                     -- width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal width_adapter_002_src_data                                                                          : std_logic_vector(79 downto 0); -- width_adapter_002:out_data -> burst_adapter_001:sink0_data
	signal width_adapter_002_src_ready                                                                         : std_logic;                     -- burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                       : std_logic_vector(22 downto 0); -- width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	signal id_router_021_src_endofpacket                                                                       : std_logic;                     -- id_router_021:src_endofpacket -> width_adapter_003:in_endofpacket
	signal id_router_021_src_valid                                                                             : std_logic;                     -- id_router_021:src_valid -> width_adapter_003:in_valid
	signal id_router_021_src_startofpacket                                                                     : std_logic;                     -- id_router_021:src_startofpacket -> width_adapter_003:in_startofpacket
	signal id_router_021_src_data                                                                              : std_logic_vector(79 downto 0); -- id_router_021:src_data -> width_adapter_003:in_data
	signal id_router_021_src_channel                                                                           : std_logic_vector(22 downto 0); -- id_router_021:src_channel -> width_adapter_003:in_channel
	signal id_router_021_src_ready                                                                             : std_logic;                     -- width_adapter_003:in_ready -> id_router_021:src_ready
	signal width_adapter_003_src_endofpacket                                                                   : std_logic;                     -- width_adapter_003:out_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	signal width_adapter_003_src_valid                                                                         : std_logic;                     -- width_adapter_003:out_valid -> rsp_xbar_demux_021:sink_valid
	signal width_adapter_003_src_startofpacket                                                                 : std_logic;                     -- width_adapter_003:out_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	signal width_adapter_003_src_data                                                                          : std_logic_vector(97 downto 0); -- width_adapter_003:out_data -> rsp_xbar_demux_021:sink_data
	signal width_adapter_003_src_ready                                                                         : std_logic;                     -- rsp_xbar_demux_021:sink_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                       : std_logic_vector(22 downto 0); -- width_adapter_003:out_channel -> rsp_xbar_demux_021:sink_channel
	signal limiter_cmd_valid_data                                                                              : std_logic_vector(22 downto 0); -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal limiter_001_cmd_valid_data                                                                          : std_logic_vector(22 downto 0); -- limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	signal irq_mapper_receiver0_irq                                                                            : std_logic;                     -- timer_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                            : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                            : std_logic;                     -- kb_irq:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                                            : std_logic;                     -- kick_irq:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                                            : std_logic;                     -- snare_irq:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                                            : std_logic;                     -- hh_irq:irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                                                            : std_logic;                     -- clap_irq:irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                                                            : std_logic;                     -- dac_irq:irq -> irq_mapper:receiver7_irq
	signal irq_mapper_receiver8_irq                                                                            : std_logic;                     -- timer_1:irq -> irq_mapper:receiver8_irq
	signal nios2_qsys_0_d_irq_irq                                                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	signal reset_100_reset_n_ports_inv                                                                         : std_logic;                     -- reset_100_reset_n:inv -> rst_controller:reset_in1
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                        : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart_0:av_write_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                         : std_logic;                     -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart_0:av_read_n
	signal audio_sos_s1_translator_avalon_anti_slave_0_write_ports_inv                                         : std_logic;                     -- audio_sos_s1_translator_avalon_anti_slave_0_write:inv -> audio_sos:write_n
	signal dac_irq_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                     -- dac_irq_s1_translator_avalon_anti_slave_0_write:inv -> dac_irq:write_n
	signal clap_irq_s1_translator_avalon_anti_slave_0_write_ports_inv                                          : std_logic;                     -- clap_irq_s1_translator_avalon_anti_slave_0_write:inv -> clap_irq:write_n
	signal hh_irq_s1_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                     -- hh_irq_s1_translator_avalon_anti_slave_0_write:inv -> hh_irq:write_n
	signal snare_irq_s1_translator_avalon_anti_slave_0_write_ports_inv                                         : std_logic;                     -- snare_irq_s1_translator_avalon_anti_slave_0_write:inv -> snare_irq:write_n
	signal kick_irq_s1_translator_avalon_anti_slave_0_write_ports_inv                                          : std_logic;                     -- kick_irq_s1_translator_avalon_anti_slave_0_write:inv -> kick_irq:write_n
	signal kb_irq_s1_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                     -- kb_irq_s1_translator_avalon_anti_slave_0_write:inv -> kb_irq:write_n
	signal seq_hh_s1_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                     -- seq_hh_s1_translator_avalon_anti_slave_0_write:inv -> seq_hh:write_n
	signal seq_snare_s1_translator_avalon_anti_slave_0_write_ports_inv                                         : std_logic;                     -- seq_snare_s1_translator_avalon_anti_slave_0_write:inv -> seq_snare:write_n
	signal led_r_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                     -- led_r_s1_translator_avalon_anti_slave_0_write:inv -> led_r:write_n
	signal timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                     -- timer_0_s1_translator_avalon_anti_slave_0_write:inv -> timer_0:write_n
	signal seq_clap_s1_translator_avalon_anti_slave_0_write_ports_inv                                          : std_logic;                     -- seq_clap_s1_translator_avalon_anti_slave_0_write:inv -> seq_clap:write_n
	signal seq_kick_s1_translator_avalon_anti_slave_0_write_ports_inv                                          : std_logic;                     -- seq_kick_s1_translator_avalon_anti_slave_0_write:inv -> seq_kick:write_n
	signal wr_address_s1_translator_avalon_anti_slave_0_write_ports_inv                                        : std_logic;                     -- wr_address_s1_translator_avalon_anti_slave_0_write:inv -> wr_address:write_n
	signal color_out_s1_translator_avalon_anti_slave_0_write_ports_inv                                         : std_logic;                     -- color_out_s1_translator_avalon_anti_slave_0_write:inv -> color_out:write_n
	signal wr_en_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                     -- wr_en_s1_translator_avalon_anti_slave_0_write:inv -> wr_en:write_n
	signal timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                     -- timer_1_s1_translator_avalon_anti_slave_0_write:inv -> timer_1:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [AUDIO_DAC_FIFO_0:reset_n, SRAM_DE2_0:reset_n, audio_sos:reset_n, clap_irq:reset_n, color_out:reset_n, dac_irq:reset_n, hh_irq:reset_n, in_bus:reset_n, jtag_uart_0:rst_n, kb_data:reset_n, kb_irq:reset_n, kick_irq:reset_n, led_r:reset_n, nios2_qsys_0:reset_n, seq_clap:reset_n, seq_hh:reset_n, seq_kick:reset_n, seq_snare:reset_n, snare_irq:reset_n, timer_0:reset_n, timer_1:reset_n, wr_address:reset_n, wr_en:reset_n]

begin

	sram_de2_0 : component SRAM_DE2
		port map (
			clk               => clk_100_clk,                                             --         clock.clk
			reset_n           => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			avs_s0_readdata   => sram_de2_0_s0_translator_avalon_anti_slave_0_readdata,   --            s0.readdata
			avs_s0_writedata  => sram_de2_0_s0_translator_avalon_anti_slave_0_writedata,  --              .writedata
			avs_s0_address    => sram_de2_0_s0_translator_avalon_anti_slave_0_address,    --              .address
			avs_s0_write      => sram_de2_0_s0_translator_avalon_anti_slave_0_write,      --              .write
			avs_s0_read       => sram_de2_0_s0_translator_avalon_anti_slave_0_read,       --              .read
			avs_s0_byteenable => sram_de2_0_s0_translator_avalon_anti_slave_0_byteenable, --              .byteenable
			coe_SRAM_ADDR     => sram_de2_ADDR,                                           -- conduit_end_0.export
			coe_SRAM_DQ       => sram_de2_DQ,                                             --              .export
			coe_SRAM_WE_N     => sram_de2_WE_N,                                           --              .export
			coe_SRAM_OE_N     => sram_de2_OE_N,                                           --              .export
			coe_SRAM_UB_N     => sram_de2_UB_N,                                           --              .export
			coe_SRAM_LB_N     => sram_de2_LB_N,                                           --              .export
			coe_SRAM_CE_N     => sram_de2_CE_N                                            --              .export
		);

	nios2_qsys_0 : component nios_ii_nios2_qsys_0
		port map (
			clk                                   => clk_100_clk,                                                               --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                                  --                   reset_n.reset_n
			d_address                             => nios2_qsys_0_data_master_address,                                          --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                                       --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                             --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                                            --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                                        --                          .writedata
			d_readdatavalid                       => nios2_qsys_0_data_master_readdatavalid,                                    --                          .readdatavalid
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                                   --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                                      --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                               --                          .waitrequest
			i_readdatavalid                       => nios2_qsys_0_instruction_master_readdatavalid,                             --                          .readdatavalid
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => nios2_qsys_0_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                                       -- custom_instruction_master.readra
		);

	in_bus : component nios_ii_in_bus
		port map (
			clk      => clk_100_clk,                                       --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address  => in_bus_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => in_bus_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => in_bus_export                                      -- external_connection.export
		);

	wr_en : component nios_ii_wr_en
		port map (
			clk        => clk_100_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => wr_en_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => wr_en_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => wr_en_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => wr_en_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => wr_en_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => wr_en_export                                             -- external_connection.export
		);

	color_out : component nios_ii_color_out
		port map (
			clk        => clk_100_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => color_out_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => color_out_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => color_out_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => color_out_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => color_out_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => color_out_export                                             -- external_connection.export
		);

	wr_address : component nios_ii_wr_address
		port map (
			clk        => clk_100_clk,                                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                     --               reset.reset_n
			address    => wr_address_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => wr_address_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => wr_address_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => wr_address_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => wr_address_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => wr_address_export                                             -- external_connection.export
		);

	seq_clap : component nios_ii_seq_clap
		port map (
			clk        => clk_100_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => seq_clap_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => seq_clap_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => seq_clap_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => seq_clap_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => seq_clap_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => seq_clap_export                                             -- external_connection.export
		);

	seq_kick : component nios_ii_seq_clap
		port map (
			clk        => clk_100_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => seq_kick_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => seq_kick_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => seq_kick_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => seq_kick_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => seq_kick_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => seq_kick_export                                             -- external_connection.export
		);

	timer_0 : component nios_ii_timer_0
		port map (
			clk        => clk_100_clk,                                               --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_0_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_0_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_0_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_0_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                                   --   irq.irq
		);

	jtag_uart_0 : component nios_ii_jtag_uart_0
		port map (
			clk            => clk_100_clk,                                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                     --             reset.reset_n
			av_chipselect  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                                      --               irq.irq
		);

	led_r : component nios_ii_led_r
		port map (
			clk        => clk_100_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => led_r_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => led_r_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => led_r_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => led_r_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => led_r_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => led_r_export                                             -- external_connection.export
		);

	seq_snare : component nios_ii_seq_clap
		port map (
			clk        => clk_100_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => seq_snare_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => seq_snare_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => seq_snare_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => seq_snare_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => seq_snare_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => seq_snare_export                                             -- external_connection.export
		);

	seq_hh : component nios_ii_seq_clap
		port map (
			clk        => clk_100_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                 --               reset.reset_n
			address    => seq_hh_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => seq_hh_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => seq_hh_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => seq_hh_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => seq_hh_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => seq_hh_export                                             -- external_connection.export
		);

	kb_irq : component nios_ii_kb_irq
		port map (
			clk        => clk_100_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                 --               reset.reset_n
			address    => kb_irq_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => kb_irq_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => kb_irq_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => kb_irq_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => kb_irq_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => kb_irq_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver2_irq                                  --                 irq.irq
		);

	kb_data : component nios_ii_kb_data
		port map (
			clk      => clk_100_clk,                                        --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,           --               reset.reset_n
			address  => kb_data_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => kb_data_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => kb_data_export                                      -- external_connection.export
		);

	kick_irq : component nios_ii_kb_irq
		port map (
			clk        => clk_100_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => kick_irq_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => kick_irq_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => kick_irq_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => kick_irq_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => kick_irq_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => kick_irq_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver3_irq                                    --                 irq.irq
		);

	snare_irq : component nios_ii_kb_irq
		port map (
			clk        => clk_100_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => snare_irq_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => snare_irq_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => snare_irq_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => snare_irq_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => snare_irq_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => snare_irq_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver4_irq                                     --                 irq.irq
		);

	hh_irq : component nios_ii_kb_irq
		port map (
			clk        => clk_100_clk,                                              --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                 --               reset.reset_n
			address    => hh_irq_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => hh_irq_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => hh_irq_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => hh_irq_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => hh_irq_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => hh_irq_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver5_irq                                  --                 irq.irq
		);

	clap_irq : component nios_ii_kb_irq
		port map (
			clk        => clk_100_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => clap_irq_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => clap_irq_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => clap_irq_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => clap_irq_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => clap_irq_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => clap_irq_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver6_irq                                    --                 irq.irq
		);

	dac_irq : component nios_ii_kb_irq
		port map (
			clk        => clk_100_clk,                                               --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  --               reset.reset_n
			address    => dac_irq_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => dac_irq_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => dac_irq_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => dac_irq_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => dac_irq_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => dac_irq_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver7_irq                                   --                 irq.irq
		);

	audio_dac_fifo_0 : component AUDIO_DAC_FIFO
		generic map (
			REF_CLK     => 18432000,
			SAMPLE_RATE => 48000,
			DATA_WIDTH  => 16,
			CHANNEL_NUM => 2
		)
		port map (
			avs_s0_writedata => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_writedata, --          s0.writedata
			avs_s0_write     => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_write,     --            .write
			avs_s0_readdata  => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_readdata,  --            .readdata
			avs_s0_read      => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_read,      --            .read
			clk              => clk_100_clk,                                                  --       clock.clk
			reset_n          => rst_controller_reset_out_reset_ports_inv,                     --       reset.reset_n
			oAUD_BCK         => audio_dac_fifo_oAUD_BCK,                                      -- conduit_end.export
			oAUD_LRCK        => audio_dac_fifo_oAUD_LRCK,                                     --            .export
			oAUD_DATA        => audio_dac_fifo_oAUD_DATA,                                     --            .export
			oAUD_XCK         => audio_dac_fifo_oAUD_XCK,                                      --            .export
			iCLK_18_4        => audio_dac_fifo_iCLK_18_4                                      --            .export
		);

	audio_sos : component nios_ii_seq_clap
		port map (
			clk        => clk_100_clk,                                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                    --               reset.reset_n
			address    => audio_sos_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => audio_sos_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => audio_sos_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => audio_sos_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => audio_sos_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => audio_sos_export                                             -- external_connection.export
		);

	timer_1 : component nios_ii_timer_0
		port map (
			clk        => clk_100_clk,                                               --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_1_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_1_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_1_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_1_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver8_irq                                   --   irq.irq
		);

	nios2_qsys_0_instruction_master_translator : component nios_ii_nios2_qsys_0_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 21,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 21,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_100_clk,                                                                        --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                                     --                     reset.reset
			uav_address              => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_qsys_0_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_qsys_0_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => nios2_qsys_0_instruction_master_read,                                               --                          .read
			av_readdata              => nios2_qsys_0_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid         => nios2_qsys_0_instruction_master_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                                --               (terminated)
			av_byteenable            => "1111",                                                                             --               (terminated)
			av_beginbursttransfer    => '0',                                                                                --               (terminated)
			av_begintransfer         => '0',                                                                                --               (terminated)
			av_chipselect            => '0',                                                                                --               (terminated)
			av_write                 => '0',                                                                                --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                                 --               (terminated)
			av_lock                  => '0',                                                                                --               (terminated)
			av_debugaccess           => '0',                                                                                --               (terminated)
			uav_clken                => open,                                                                               --               (terminated)
			av_clken                 => '1',                                                                                --               (terminated)
			uav_response             => "00",                                                                               --               (terminated)
			av_response              => open,                                                                               --               (terminated)
			uav_writeresponserequest => open,                                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                                --               (terminated)
		);

	nios2_qsys_0_data_master_translator : component nios_ii_nios2_qsys_0_data_master_translator
		generic map (
			AV_ADDRESS_W                => 21,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 21,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_100_clk,                                                                 --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                     reset.reset
			uav_address              => nios2_qsys_0_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => nios2_qsys_0_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => nios2_qsys_0_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => nios2_qsys_0_data_master_byteenable,                                         --                          .byteenable
			av_read                  => nios2_qsys_0_data_master_read,                                               --                          .read
			av_readdata              => nios2_qsys_0_data_master_readdata,                                           --                          .readdata
			av_readdatavalid         => nios2_qsys_0_data_master_readdatavalid,                                      --                          .readdatavalid
			av_write                 => nios2_qsys_0_data_master_write,                                              --                          .write
			av_writedata             => nios2_qsys_0_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => nios2_qsys_0_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                         --               (terminated)
			av_beginbursttransfer    => '0',                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                         --               (terminated)
			av_chipselect            => '0',                                                                         --               (terminated)
			av_lock                  => '0',                                                                         --               (terminated)
			uav_clken                => open,                                                                        --               (terminated)
			av_clken                 => '1',                                                                         --               (terminated)
			uav_response             => "00",                                                                        --               (terminated)
			av_response              => open,                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                         --               (terminated)
		);

	nios2_qsys_0_jtag_debug_module_translator : component nios_ii_nios2_qsys_0_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                            --                    reset.reset
			uav_address              => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                                      --              (terminated)
			av_burstcount            => open,                                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                                      --              (terminated)
			av_lock                  => open,                                                                                      --              (terminated)
			av_chipselect            => open,                                                                                      --              (terminated)
			av_clken                 => open,                                                                                      --              (terminated)
			uav_clken                => '0',                                                                                       --              (terminated)
			av_outputenable          => open,                                                                                      --              (terminated)
			uav_response             => open,                                                                                      --              (terminated)
			av_response              => "00",                                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                                        --              (terminated)
		);

	sram_de2_0_s0_translator : component nios_ii_sram_de2_0_s0_translator
		generic map (
			AV_ADDRESS_W                   => 18,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 2,
			AV_WRITE_WAIT_CYCLES           => 2,
			AV_SETUP_WAIT_CYCLES           => 2,
			AV_DATA_HOLD_CYCLES            => 2
		)
		port map (
			clk                      => clk_100_clk,                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address              => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sram_de2_0_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sram_de2_0_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sram_de2_0_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sram_de2_0_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sram_de2_0_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sram_de2_0_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_chipselect            => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator : component nios_ii_jtag_uart_0_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                           --                    reset.reset
			uav_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                                     --              (terminated)
			av_burstcount            => open,                                                                                     --              (terminated)
			av_byteenable            => open,                                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                                     --              (terminated)
			av_lock                  => open,                                                                                     --              (terminated)
			av_clken                 => open,                                                                                     --              (terminated)
			uav_clken                => '0',                                                                                      --              (terminated)
			av_debugaccess           => open,                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                     --              (terminated)
			uav_response             => open,                                                                                     --              (terminated)
			av_response              => "00",                                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                                       --              (terminated)
		);

	audio_sos_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => audio_sos_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => audio_sos_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => audio_sos_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => audio_sos_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => audio_sos_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	dac_irq_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => dac_irq_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => dac_irq_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => dac_irq_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => dac_irq_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => dac_irq_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	clap_irq_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address              => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => clap_irq_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => clap_irq_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => clap_irq_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => clap_irq_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => clap_irq_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	hh_irq_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => hh_irq_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => hh_irq_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => hh_irq_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => hh_irq_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => hh_irq_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	snare_irq_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => snare_irq_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => snare_irq_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => snare_irq_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => snare_irq_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => snare_irq_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	kick_irq_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address              => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => kick_irq_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => kick_irq_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => kick_irq_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => kick_irq_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => kick_irq_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	kb_irq_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => kb_irq_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => kb_irq_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => kb_irq_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => kb_irq_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => kb_irq_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	seq_hh_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => seq_hh_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => seq_hh_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => seq_hh_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => seq_hh_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => seq_hh_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	seq_snare_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => seq_snare_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => seq_snare_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => seq_snare_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => seq_snare_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => seq_snare_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	led_r_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => led_r_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => led_r_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => led_r_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => led_r_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => led_r_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => led_r_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => led_r_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => led_r_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => led_r_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => led_r_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => led_r_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => led_r_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => led_r_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => led_r_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => led_r_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => led_r_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                --              (terminated)
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_byteenable            => open,                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                 --              (terminated)
			av_waitrequest           => '0',                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	timer_0_s1_translator : component nios_ii_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	seq_clap_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address              => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => seq_clap_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => seq_clap_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => seq_clap_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => seq_clap_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => seq_clap_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	seq_kick_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address              => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => seq_kick_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => seq_kick_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => seq_kick_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => seq_kick_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => seq_kick_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	wr_address_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address              => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => wr_address_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => wr_address_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => wr_address_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => wr_address_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => wr_address_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	color_out_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                             --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => color_out_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => color_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => color_out_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => color_out_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => color_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => color_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => color_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => color_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => color_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => color_out_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => color_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => color_out_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => color_out_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => color_out_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => color_out_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => color_out_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	in_bus_s1_translator : component nios_ii_in_bus_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                          --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => in_bus_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => in_bus_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                 --              (terminated)
			av_read                  => open,                                                                 --              (terminated)
			av_writedata             => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_chipselect            => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	wr_en_s1_translator : component nios_ii_audio_sos_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                         --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                    reset.reset
			uav_address              => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => wr_en_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => wr_en_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => wr_en_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => wr_en_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => wr_en_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                --              (terminated)
			av_begintransfer         => open,                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                --              (terminated)
			av_burstcount            => open,                                                                --              (terminated)
			av_byteenable            => open,                                                                --              (terminated)
			av_readdatavalid         => '0',                                                                 --              (terminated)
			av_waitrequest           => '0',                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                --              (terminated)
			av_lock                  => open,                                                                --              (terminated)
			av_clken                 => open,                                                                --              (terminated)
			uav_clken                => '0',                                                                 --              (terminated)
			av_debugaccess           => open,                                                                --              (terminated)
			av_outputenable          => open,                                                                --              (terminated)
			uav_response             => open,                                                                --              (terminated)
			av_response              => "00",                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                  --              (terminated)
		);

	kb_data_s1_translator : component nios_ii_in_bus_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => kb_data_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => kb_data_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                  --              (terminated)
			av_read                  => open,                                                                  --              (terminated)
			av_writedata             => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_chipselect            => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	audio_dac_fifo_0_s0_translator : component nios_ii_audio_dac_fifo_0_s0_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                                    --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address              => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_write                 => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_write,                       --      avalon_anti_slave_0.write
			av_read                  => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => audio_dac_fifo_0_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_address               => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	timer_1_s1_translator : component nios_ii_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 21,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_100_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_1_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_1_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_1_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_BEGIN_BURST           => 76,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			PKT_BURST_TYPE_H          => 73,
			PKT_BURST_TYPE_L          => 72,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_TRANS_EXCLUSIVE       => 62,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_THREAD_ID_H           => 88,
			PKT_THREAD_ID_L           => 88,
			PKT_CACHE_H               => 95,
			PKT_CACHE_L               => 92,
			PKT_DATA_SIDEBAND_H       => 75,
			PKT_DATA_SIDEBAND_L       => 75,
			PKT_QOS_H                 => 77,
			PKT_QOS_L                 => 77,
			PKT_ADDR_SIDEBAND_H       => 74,
			PKT_ADDR_SIDEBAND_L       => 74,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			ST_DATA_W                 => 98,
			ST_CHANNEL_W              => 23,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                                 --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			av_address              => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_rsp_src_valid,                                                                       --        rp.valid
			rp_data                 => limiter_rsp_src_data,                                                                        --          .data
			rp_channel              => limiter_rsp_src_channel,                                                                     --          .channel
			rp_startofpacket        => limiter_rsp_src_startofpacket,                                                               --          .startofpacket
			rp_endofpacket          => limiter_rsp_src_endofpacket,                                                                 --          .endofpacket
			rp_ready                => limiter_rsp_src_ready,                                                                       --          .ready
			av_response             => open,                                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                                         -- (terminated)
		);

	nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_BEGIN_BURST           => 76,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			PKT_BURST_TYPE_H          => 73,
			PKT_BURST_TYPE_L          => 72,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_TRANS_EXCLUSIVE       => 62,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_THREAD_ID_H           => 88,
			PKT_THREAD_ID_L           => 88,
			PKT_CACHE_H               => 95,
			PKT_CACHE_L               => 92,
			PKT_DATA_SIDEBAND_H       => 75,
			PKT_DATA_SIDEBAND_L       => 75,
			PKT_QOS_H                 => 77,
			PKT_QOS_L                 => 77,
			PKT_ADDR_SIDEBAND_H       => 74,
			PKT_ADDR_SIDEBAND_L       => 74,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			ST_DATA_W                 => 98,
			ST_CHANNEL_W              => 23,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                          --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			av_address              => nios2_qsys_0_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_001_rsp_src_valid,                                                            --        rp.valid
			rp_data                 => limiter_001_rsp_src_data,                                                             --          .data
			rp_channel              => limiter_001_rsp_src_channel,                                                          --          .channel
			rp_startofpacket        => limiter_001_rsp_src_startofpacket,                                                    --          .startofpacket
			rp_endofpacket          => limiter_001_rsp_src_endofpacket,                                                      --          .endofpacket
			rp_ready                => limiter_001_rsp_src_ready,                                                            --          .ready
			av_response             => open,                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                  -- (terminated)
		);

	nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                      --       clk_reset.reset
			m0_address              => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                              --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                              --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                               --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                        --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                            --                .channel
			rf_sink_ready           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                  --     (terminated)
		);

	nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                      -- clk_reset.reset
			in_data           => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                -- (terminated)
			csr_read          => '0',                                                                                                 -- (terminated)
			csr_write         => '0',                                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                  -- (terminated)
			almost_full_data  => open,                                                                                                -- (terminated)
			almost_empty_data => open,                                                                                                -- (terminated)
			in_empty          => '0',                                                                                                 -- (terminated)
			out_empty         => open,                                                                                                -- (terminated)
			in_error          => '0',                                                                                                 -- (terminated)
			out_error         => open,                                                                                                -- (terminated)
			in_channel        => '0',                                                                                                 -- (terminated)
			out_channel       => open                                                                                                 -- (terminated)
		);

	sram_de2_0_s0_translator_avalon_universal_slave_0_agent : component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 58,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 38,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 39,
			PKT_TRANS_POSTED          => 40,
			PKT_TRANS_WRITE           => 41,
			PKT_TRANS_READ            => 42,
			PKT_TRANS_LOCK            => 43,
			PKT_SRC_ID_H              => 64,
			PKT_SRC_ID_L              => 60,
			PKT_DEST_ID_H             => 69,
			PKT_DEST_ID_L             => 65,
			PKT_BURSTWRAP_H           => 50,
			PKT_BURSTWRAP_L           => 48,
			PKT_BYTE_CNT_H            => 47,
			PKT_BYTE_CNT_L            => 45,
			PKT_PROTECTION_H          => 73,
			PKT_PROTECTION_L          => 71,
			PKT_RESPONSE_STATUS_H     => 79,
			PKT_RESPONSE_STATUS_L     => 78,
			PKT_BURST_SIZE_H          => 53,
			PKT_BURST_SIZE_L          => 51,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 80,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                        --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                        --                .valid
			cp_data                 => burst_adapter_source0_data,                                                         --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                  --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                      --                .channel
			rf_sink_ready           => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 81,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_002_src_ready,                                                                         --              cp.ready
			cp_valid                => cmd_xbar_mux_002_src_valid,                                                                         --                .valid
			cp_data                 => cmd_xbar_mux_002_src_data,                                                                          --                .data
			cp_startofpacket        => cmd_xbar_mux_002_src_startofpacket,                                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_002_src_endofpacket,                                                                   --                .endofpacket
			cp_channel              => cmd_xbar_mux_002_src_channel,                                                                       --                .channel
			rf_sink_ready           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                 --     (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                               -- (terminated)
			csr_read          => '0',                                                                                                -- (terminated)
			csr_write         => '0',                                                                                                -- (terminated)
			csr_readdata      => open,                                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                 -- (terminated)
			almost_full_data  => open,                                                                                               -- (terminated)
			almost_empty_data => open,                                                                                               -- (terminated)
			in_empty          => '0',                                                                                                -- (terminated)
			out_empty         => open,                                                                                               -- (terminated)
			in_error          => '0',                                                                                                -- (terminated)
			out_error         => open,                                                                                               -- (terminated)
			in_channel        => '0',                                                                                                -- (terminated)
			out_channel       => open                                                                                                -- (terminated)
		);

	audio_sos_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => audio_sos_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_003_src_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_mux_003_src_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_mux_003_src_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_mux_003_src_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_003_src_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_mux_003_src_channel,                                                      --                .channel
			rf_sink_ready           => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => audio_sos_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => audio_sos_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => audio_sos_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	dac_irq_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => dac_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_004_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_004_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_004_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_004_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_004_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_004_src_channel,                                                    --                .channel
			rf_sink_ready           => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => dac_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => dac_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => dac_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	clap_irq_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => clap_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_005_src_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_mux_005_src_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_mux_005_src_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_mux_005_src_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_005_src_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_mux_005_src_channel,                                                     --                .channel
			rf_sink_ready           => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => clap_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => clap_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => clap_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	hh_irq_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => hh_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_006_src_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_006_src_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_mux_006_src_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_006_src_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_006_src_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_006_src_channel,                                                   --                .channel
			rf_sink_ready           => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => hh_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => hh_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => hh_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	snare_irq_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => snare_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_007_src_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_mux_007_src_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_mux_007_src_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_mux_007_src_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_007_src_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_mux_007_src_channel,                                                      --                .channel
			rf_sink_ready           => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => snare_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => snare_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => snare_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	kick_irq_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => kick_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_008_src_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_mux_008_src_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_mux_008_src_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_mux_008_src_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_008_src_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_mux_008_src_channel,                                                     --                .channel
			rf_sink_ready           => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => kick_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => kick_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => kick_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	kb_irq_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => kb_irq_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_009_src_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_009_src_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_mux_009_src_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_009_src_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_009_src_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_009_src_channel,                                                   --                .channel
			rf_sink_ready           => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => kb_irq_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => kb_irq_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => kb_irq_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	seq_hh_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => seq_hh_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_010_src_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_010_src_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_mux_010_src_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_010_src_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_010_src_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_010_src_channel,                                                   --                .channel
			rf_sink_ready           => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => seq_hh_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => seq_hh_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => seq_hh_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	seq_snare_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => seq_snare_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_011_src_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_mux_011_src_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_mux_011_src_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_mux_011_src_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_011_src_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_mux_011_src_channel,                                                      --                .channel
			rf_sink_ready           => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => seq_snare_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => seq_snare_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => seq_snare_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	led_r_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => led_r_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => led_r_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => led_r_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => led_r_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => led_r_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => led_r_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => led_r_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => led_r_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => led_r_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => led_r_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => led_r_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => led_r_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => led_r_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => led_r_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => led_r_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => led_r_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_012_src_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_mux_012_src_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_mux_012_src_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_mux_012_src_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_012_src_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_mux_012_src_channel,                                                  --                .channel
			rf_sink_ready           => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => led_r_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => led_r_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => led_r_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_013_src_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_013_src_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_mux_013_src_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_013_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_013_src_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_013_src_channel,                                                    --                .channel
			rf_sink_ready           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	seq_clap_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => seq_clap_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_014_src_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_mux_014_src_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_mux_014_src_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_mux_014_src_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_014_src_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_mux_014_src_channel,                                                     --                .channel
			rf_sink_ready           => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => seq_clap_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => seq_clap_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => seq_clap_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	seq_kick_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => seq_kick_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_015_src_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_mux_015_src_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_mux_015_src_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_mux_015_src_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_015_src_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_mux_015_src_channel,                                                     --                .channel
			rf_sink_ready           => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => seq_kick_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => seq_kick_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => seq_kick_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	wr_address_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => wr_address_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_016_src_ready,                                                         --              cp.ready
			cp_valid                => cmd_xbar_mux_016_src_valid,                                                         --                .valid
			cp_data                 => cmd_xbar_mux_016_src_data,                                                          --                .data
			cp_startofpacket        => cmd_xbar_mux_016_src_startofpacket,                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_016_src_endofpacket,                                                   --                .endofpacket
			cp_channel              => cmd_xbar_mux_016_src_channel,                                                       --                .channel
			rf_sink_ready           => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => wr_address_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => wr_address_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => wr_address_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	color_out_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => color_out_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => color_out_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => color_out_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => color_out_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => color_out_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => color_out_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => color_out_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => color_out_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => color_out_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => color_out_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => color_out_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => color_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => color_out_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => color_out_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => color_out_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => color_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_017_src_ready,                                                        --              cp.ready
			cp_valid                => cmd_xbar_mux_017_src_valid,                                                        --                .valid
			cp_data                 => cmd_xbar_mux_017_src_data,                                                         --                .data
			cp_startofpacket        => cmd_xbar_mux_017_src_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_017_src_endofpacket,                                                  --                .endofpacket
			cp_channel              => cmd_xbar_mux_017_src_channel,                                                      --                .channel
			rf_sink_ready           => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => color_out_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => color_out_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => color_out_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	in_bus_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                    --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => in_bus_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_018_src_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_mux_018_src_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_mux_018_src_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_mux_018_src_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_018_src_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_mux_018_src_channel,                                                   --                .channel
			rf_sink_ready           => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => in_bus_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                    --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => in_bus_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => in_bus_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	wr_en_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                   --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => wr_en_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_019_src_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_mux_019_src_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_mux_019_src_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_mux_019_src_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_019_src_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_mux_019_src_channel,                                                  --                .channel
			rf_sink_ready           => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => wr_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                            --     (terminated)
		);

	wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			in_data           => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => wr_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => wr_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                          -- (terminated)
			csr_read          => '0',                                                                           -- (terminated)
			csr_write         => '0',                                                                           -- (terminated)
			csr_readdata      => open,                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                            -- (terminated)
			almost_full_data  => open,                                                                          -- (terminated)
			almost_empty_data => open,                                                                          -- (terminated)
			in_empty          => '0',                                                                           -- (terminated)
			out_empty         => open,                                                                          -- (terminated)
			in_error          => '0',                                                                           -- (terminated)
			out_error         => open,                                                                          -- (terminated)
			in_channel        => '0',                                                                           -- (terminated)
			out_channel       => open                                                                           -- (terminated)
		);

	kb_data_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => kb_data_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src20_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src20_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src20_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src20_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src20_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src20_channel,                                                --                .channel
			rf_sink_ready           => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => kb_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => kb_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => kb_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent : component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 58,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 38,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 39,
			PKT_TRANS_POSTED          => 40,
			PKT_TRANS_WRITE           => 41,
			PKT_TRANS_READ            => 42,
			PKT_TRANS_LOCK            => 43,
			PKT_SRC_ID_H              => 64,
			PKT_SRC_ID_L              => 60,
			PKT_DEST_ID_H             => 69,
			PKT_DEST_ID_L             => 65,
			PKT_BURSTWRAP_H           => 50,
			PKT_BURSTWRAP_L           => 48,
			PKT_BYTE_CNT_H            => 47,
			PKT_BYTE_CNT_L            => 45,
			PKT_PROTECTION_H          => 73,
			PKT_PROTECTION_L          => 71,
			PKT_RESPONSE_STATUS_H     => 79,
			PKT_RESPONSE_STATUS_L     => 78,
			PKT_BURST_SIZE_H          => 53,
			PKT_BURST_SIZE_L          => 51,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 80,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                          --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                          --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                           --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                                  --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                                    --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                        --                .channel
			rf_sink_ready           => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 81,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 56,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 57,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			PKT_TRANS_READ            => 60,
			PKT_TRANS_LOCK            => 61,
			PKT_SRC_ID_H              => 82,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 66,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_PROTECTION_H          => 91,
			PKT_PROTECTION_L          => 89,
			PKT_RESPONSE_STATUS_H     => 97,
			PKT_RESPONSE_STATUS_L     => 96,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 23,
			ST_DATA_W                 => 98,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_100_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src22_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src22_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src22_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src22_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src22_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src22_channel,                                                --                .channel
			rf_sink_ready           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component nios_ii_nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 99,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_100_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	addr_router : component nios_ii_addr_router
		port map (
			sink_ready         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                                                 --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                       --       src.ready
			src_valid          => addr_router_src_valid,                                                                       --          .valid
			src_data           => addr_router_src_data,                                                                        --          .data
			src_channel        => addr_router_src_channel,                                                                     --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                  --          .endofpacket
		);

	addr_router_001 : component nios_ii_addr_router_001
		port map (
			sink_ready         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                            --       src.ready
			src_valid          => addr_router_001_src_valid,                                                            --          .valid
			src_data           => addr_router_001_src_data,                                                             --          .data
			src_channel        => addr_router_001_src_channel,                                                          --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                       --          .endofpacket
		);

	id_router : component nios_ii_id_router
		port map (
			sink_ready         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                       --       src.ready
			src_valid          => id_router_src_valid,                                                                       --          .valid
			src_data           => id_router_src_data,                                                                        --          .data
			src_channel        => id_router_src_channel,                                                                     --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                               --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                                  --          .endofpacket
		);

	id_router_001 : component nios_ii_id_router_001
		port map (
			sink_ready         => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sram_de2_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                  --       src.ready
			src_valid          => id_router_001_src_valid,                                                  --          .valid
			src_data           => id_router_001_src_data,                                                   --          .data
			src_channel        => id_router_001_src_channel,                                                --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                             --          .endofpacket
		);

	id_router_002 : component nios_ii_id_router
		port map (
			sink_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                  --       src.ready
			src_valid          => id_router_002_src_valid,                                                                  --          .valid
			src_data           => id_router_002_src_data,                                                                   --          .data
			src_channel        => id_router_002_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                             --          .endofpacket
		);

	id_router_003 : component nios_ii_id_router
		port map (
			sink_ready         => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => audio_sos_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                 --       src.ready
			src_valid          => id_router_003_src_valid,                                                 --          .valid
			src_data           => id_router_003_src_data,                                                  --          .data
			src_channel        => id_router_003_src_channel,                                               --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                            --          .endofpacket
		);

	id_router_004 : component nios_ii_id_router
		port map (
			sink_ready         => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => dac_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                               --       src.ready
			src_valid          => id_router_004_src_valid,                                               --          .valid
			src_data           => id_router_004_src_data,                                                --          .data
			src_channel        => id_router_004_src_channel,                                             --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                          --          .endofpacket
		);

	id_router_005 : component nios_ii_id_router
		port map (
			sink_ready         => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => clap_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                --       src.ready
			src_valid          => id_router_005_src_valid,                                                --          .valid
			src_data           => id_router_005_src_data,                                                 --          .data
			src_channel        => id_router_005_src_channel,                                              --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                           --          .endofpacket
		);

	id_router_006 : component nios_ii_id_router
		port map (
			sink_ready         => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => hh_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                              --       src.ready
			src_valid          => id_router_006_src_valid,                                              --          .valid
			src_data           => id_router_006_src_data,                                               --          .data
			src_channel        => id_router_006_src_channel,                                            --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                         --          .endofpacket
		);

	id_router_007 : component nios_ii_id_router
		port map (
			sink_ready         => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => snare_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                 --       src.ready
			src_valid          => id_router_007_src_valid,                                                 --          .valid
			src_data           => id_router_007_src_data,                                                  --          .data
			src_channel        => id_router_007_src_channel,                                               --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                            --          .endofpacket
		);

	id_router_008 : component nios_ii_id_router
		port map (
			sink_ready         => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => kick_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                --       src.ready
			src_valid          => id_router_008_src_valid,                                                --          .valid
			src_data           => id_router_008_src_data,                                                 --          .data
			src_channel        => id_router_008_src_channel,                                              --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                           --          .endofpacket
		);

	id_router_009 : component nios_ii_id_router
		port map (
			sink_ready         => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => kb_irq_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                              --       src.ready
			src_valid          => id_router_009_src_valid,                                              --          .valid
			src_data           => id_router_009_src_data,                                               --          .data
			src_channel        => id_router_009_src_channel,                                            --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                         --          .endofpacket
		);

	id_router_010 : component nios_ii_id_router
		port map (
			sink_ready         => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => seq_hh_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                              --       src.ready
			src_valid          => id_router_010_src_valid,                                              --          .valid
			src_data           => id_router_010_src_data,                                               --          .data
			src_channel        => id_router_010_src_channel,                                            --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                         --          .endofpacket
		);

	id_router_011 : component nios_ii_id_router
		port map (
			sink_ready         => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => seq_snare_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                 --       src.ready
			src_valid          => id_router_011_src_valid,                                                 --          .valid
			src_data           => id_router_011_src_data,                                                  --          .data
			src_channel        => id_router_011_src_channel,                                               --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                            --          .endofpacket
		);

	id_router_012 : component nios_ii_id_router
		port map (
			sink_ready         => led_r_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => led_r_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => led_r_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => led_r_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => led_r_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                             --       src.ready
			src_valid          => id_router_012_src_valid,                                             --          .valid
			src_data           => id_router_012_src_data,                                              --          .data
			src_channel        => id_router_012_src_channel,                                           --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                        --          .endofpacket
		);

	id_router_013 : component nios_ii_id_router
		port map (
			sink_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                               --       src.ready
			src_valid          => id_router_013_src_valid,                                               --          .valid
			src_data           => id_router_013_src_data,                                                --          .data
			src_channel        => id_router_013_src_channel,                                             --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                          --          .endofpacket
		);

	id_router_014 : component nios_ii_id_router
		port map (
			sink_ready         => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => seq_clap_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                                --       src.ready
			src_valid          => id_router_014_src_valid,                                                --          .valid
			src_data           => id_router_014_src_data,                                                 --          .data
			src_channel        => id_router_014_src_channel,                                              --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                           --          .endofpacket
		);

	id_router_015 : component nios_ii_id_router
		port map (
			sink_ready         => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => seq_kick_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_015_src_ready,                                                --       src.ready
			src_valid          => id_router_015_src_valid,                                                --          .valid
			src_data           => id_router_015_src_data,                                                 --          .data
			src_channel        => id_router_015_src_channel,                                              --          .channel
			src_startofpacket  => id_router_015_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_015_src_endofpacket                                           --          .endofpacket
		);

	id_router_016 : component nios_ii_id_router
		port map (
			sink_ready         => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => wr_address_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_016_src_ready,                                                  --       src.ready
			src_valid          => id_router_016_src_valid,                                                  --          .valid
			src_data           => id_router_016_src_data,                                                   --          .data
			src_channel        => id_router_016_src_channel,                                                --          .channel
			src_startofpacket  => id_router_016_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_016_src_endofpacket                                             --          .endofpacket
		);

	id_router_017 : component nios_ii_id_router
		port map (
			sink_ready         => color_out_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => color_out_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => color_out_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => color_out_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => color_out_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_017_src_ready,                                                 --       src.ready
			src_valid          => id_router_017_src_valid,                                                 --          .valid
			src_data           => id_router_017_src_data,                                                  --          .data
			src_channel        => id_router_017_src_channel,                                               --          .channel
			src_startofpacket  => id_router_017_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_017_src_endofpacket                                            --          .endofpacket
		);

	id_router_018 : component nios_ii_id_router
		port map (
			sink_ready         => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => in_bus_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                          --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_018_src_ready,                                              --       src.ready
			src_valid          => id_router_018_src_valid,                                              --          .valid
			src_data           => id_router_018_src_data,                                               --          .data
			src_channel        => id_router_018_src_channel,                                            --          .channel
			src_startofpacket  => id_router_018_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_018_src_endofpacket                                         --          .endofpacket
		);

	id_router_019 : component nios_ii_id_router
		port map (
			sink_ready         => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => wr_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                         --       clk.clk
			reset              => rst_controller_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_019_src_ready,                                             --       src.ready
			src_valid          => id_router_019_src_valid,                                             --          .valid
			src_data           => id_router_019_src_data,                                              --          .data
			src_channel        => id_router_019_src_channel,                                           --          .channel
			src_startofpacket  => id_router_019_src_startofpacket,                                     --          .startofpacket
			src_endofpacket    => id_router_019_src_endofpacket                                        --          .endofpacket
		);

	id_router_020 : component nios_ii_id_router_020
		port map (
			sink_ready         => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => kb_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_020_src_ready,                                               --       src.ready
			src_valid          => id_router_020_src_valid,                                               --          .valid
			src_data           => id_router_020_src_data,                                                --          .data
			src_channel        => id_router_020_src_channel,                                             --          .channel
			src_startofpacket  => id_router_020_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_020_src_endofpacket                                          --          .endofpacket
		);

	id_router_021 : component nios_ii_id_router_021
		port map (
			sink_ready         => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => audio_dac_fifo_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_021_src_ready,                                                        --       src.ready
			src_valid          => id_router_021_src_valid,                                                        --          .valid
			src_data           => id_router_021_src_data,                                                         --          .data
			src_channel        => id_router_021_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_021_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_021_src_endofpacket                                                   --          .endofpacket
		);

	id_router_022 : component nios_ii_id_router_020
		port map (
			sink_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_100_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_022_src_ready,                                               --       src.ready
			src_valid          => id_router_022_src_valid,                                               --          .valid
			src_data           => id_router_022_src_data,                                                --          .data
			src_channel        => id_router_022_src_channel,                                             --          .channel
			src_startofpacket  => id_router_022_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_022_src_endofpacket                                          --          .endofpacket
		);

	limiter : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			MAX_OUTSTANDING_RESPONSES => 3,
			PIPELINED                 => 0,
			ST_DATA_W                 => 98,
			ST_CHANNEL_W              => 23,
			VALID_WIDTH               => 23,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_100_clk,                    --       clk.clk
			reset                  => rst_controller_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,          --          .valid
			cmd_sink_data          => addr_router_src_data,           --          .data
			cmd_sink_channel       => addr_router_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data          -- cmd_valid.data
		);

	limiter_001 : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 87,
			PKT_DEST_ID_L             => 83,
			PKT_TRANS_POSTED          => 58,
			PKT_TRANS_WRITE           => 59,
			MAX_OUTSTANDING_RESPONSES => 3,
			PIPELINED                 => 0,
			ST_DATA_W                 => 98,
			ST_CHANNEL_W              => 23,
			VALID_WIDTH               => 23,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 65,
			PKT_BYTE_CNT_L            => 63,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_100_clk,                        --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_001_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_001_src_valid,          --          .valid
			cmd_sink_data          => addr_router_001_src_data,           --          .data
			cmd_sink_channel       => addr_router_001_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_001_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_001_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_001_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_001_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_001_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_001_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_001_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_001_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_001_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_001_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_001_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_001_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_001_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_001_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_001_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_001_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_001_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_001_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_001_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_001_cmd_valid_data          -- cmd_valid.data
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 38,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 58,
			PKT_BYTE_CNT_H            => 47,
			PKT_BYTE_CNT_L            => 45,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 53,
			PKT_BURST_SIZE_L          => 51,
			PKT_BURST_TYPE_H          => 55,
			PKT_BURST_TYPE_L          => 54,
			PKT_BURSTWRAP_H           => 50,
			PKT_BURSTWRAP_L           => 48,
			PKT_TRANS_COMPRESSED_READ => 39,
			PKT_TRANS_WRITE           => 41,
			PKT_TRANS_READ            => 42,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 80,
			ST_CHANNEL_W              => 23,
			OUT_BYTE_CNT_H            => 46,
			OUT_BURSTWRAP_H           => 50,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => clk_100_clk,                         --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 38,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 58,
			PKT_BYTE_CNT_H            => 47,
			PKT_BYTE_CNT_L            => 45,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 53,
			PKT_BURST_SIZE_L          => 51,
			PKT_BURST_TYPE_H          => 55,
			PKT_BURST_TYPE_L          => 54,
			PKT_BURSTWRAP_H           => 50,
			PKT_BURSTWRAP_L           => 48,
			PKT_TRANS_COMPRESSED_READ => 39,
			PKT_TRANS_WRITE           => 41,
			PKT_TRANS_READ            => 42,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 80,
			ST_CHANNEL_W              => 23,
			OUT_BYTE_CNT_H            => 46,
			OUT_BURSTWRAP_H           => 50,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 7,
			BURSTWRAP_CONST_VALUE     => 7
		)
		port map (
			clk                   => clk_100_clk,                             --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => width_adapter_002_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_002_src_data,              --          .data
			sink0_channel         => width_adapter_002_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_002_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_002_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_002_src_ready,             --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2
		)
		port map (
			reset_in0  => nios2_qsys_0_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1  => reset_100_reset_n_ports_inv,                -- reset_in1.reset
			clk        => clk_100_clk,                                --       clk.clk
			reset_out  => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_in2  => '0',                                        -- (terminated)
			reset_in3  => '0',                                        -- (terminated)
			reset_in4  => '0',                                        -- (terminated)
			reset_in5  => '0',                                        -- (terminated)
			reset_in6  => '0',                                        -- (terminated)
			reset_in7  => '0',                                        -- (terminated)
			reset_in8  => '0',                                        -- (terminated)
			reset_in9  => '0',                                        -- (terminated)
			reset_in10 => '0',                                        -- (terminated)
			reset_in11 => '0',                                        -- (terminated)
			reset_in12 => '0',                                        -- (terminated)
			reset_in13 => '0',                                        -- (terminated)
			reset_in14 => '0',                                        -- (terminated)
			reset_in15 => '0'                                         -- (terminated)
		);

	cmd_xbar_demux : component nios_ii_cmd_xbar_demux
		port map (
			clk                 => clk_100_clk,                        --        clk.clk
			reset               => rst_controller_reset_out_reset,     --  clk_reset.reset
			sink_ready          => limiter_cmd_src_ready,              --       sink.ready
			sink_channel        => limiter_cmd_src_channel,            --           .channel
			sink_data           => limiter_cmd_src_data,               --           .data
			sink_startofpacket  => limiter_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket    => limiter_cmd_src_endofpacket,        --           .endofpacket
			sink_valid          => limiter_cmd_valid_data,             -- sink_valid.data
			src0_ready          => cmd_xbar_demux_src0_ready,          --       src0.ready
			src0_valid          => cmd_xbar_demux_src0_valid,          --           .valid
			src0_data           => cmd_xbar_demux_src0_data,           --           .data
			src0_channel        => cmd_xbar_demux_src0_channel,        --           .channel
			src0_startofpacket  => cmd_xbar_demux_src0_startofpacket,  --           .startofpacket
			src0_endofpacket    => cmd_xbar_demux_src0_endofpacket,    --           .endofpacket
			src1_ready          => cmd_xbar_demux_src1_ready,          --       src1.ready
			src1_valid          => cmd_xbar_demux_src1_valid,          --           .valid
			src1_data           => cmd_xbar_demux_src1_data,           --           .data
			src1_channel        => cmd_xbar_demux_src1_channel,        --           .channel
			src1_startofpacket  => cmd_xbar_demux_src1_startofpacket,  --           .startofpacket
			src1_endofpacket    => cmd_xbar_demux_src1_endofpacket,    --           .endofpacket
			src2_ready          => cmd_xbar_demux_src2_ready,          --       src2.ready
			src2_valid          => cmd_xbar_demux_src2_valid,          --           .valid
			src2_data           => cmd_xbar_demux_src2_data,           --           .data
			src2_channel        => cmd_xbar_demux_src2_channel,        --           .channel
			src2_startofpacket  => cmd_xbar_demux_src2_startofpacket,  --           .startofpacket
			src2_endofpacket    => cmd_xbar_demux_src2_endofpacket,    --           .endofpacket
			src3_ready          => cmd_xbar_demux_src3_ready,          --       src3.ready
			src3_valid          => cmd_xbar_demux_src3_valid,          --           .valid
			src3_data           => cmd_xbar_demux_src3_data,           --           .data
			src3_channel        => cmd_xbar_demux_src3_channel,        --           .channel
			src3_startofpacket  => cmd_xbar_demux_src3_startofpacket,  --           .startofpacket
			src3_endofpacket    => cmd_xbar_demux_src3_endofpacket,    --           .endofpacket
			src4_ready          => cmd_xbar_demux_src4_ready,          --       src4.ready
			src4_valid          => cmd_xbar_demux_src4_valid,          --           .valid
			src4_data           => cmd_xbar_demux_src4_data,           --           .data
			src4_channel        => cmd_xbar_demux_src4_channel,        --           .channel
			src4_startofpacket  => cmd_xbar_demux_src4_startofpacket,  --           .startofpacket
			src4_endofpacket    => cmd_xbar_demux_src4_endofpacket,    --           .endofpacket
			src5_ready          => cmd_xbar_demux_src5_ready,          --       src5.ready
			src5_valid          => cmd_xbar_demux_src5_valid,          --           .valid
			src5_data           => cmd_xbar_demux_src5_data,           --           .data
			src5_channel        => cmd_xbar_demux_src5_channel,        --           .channel
			src5_startofpacket  => cmd_xbar_demux_src5_startofpacket,  --           .startofpacket
			src5_endofpacket    => cmd_xbar_demux_src5_endofpacket,    --           .endofpacket
			src6_ready          => cmd_xbar_demux_src6_ready,          --       src6.ready
			src6_valid          => cmd_xbar_demux_src6_valid,          --           .valid
			src6_data           => cmd_xbar_demux_src6_data,           --           .data
			src6_channel        => cmd_xbar_demux_src6_channel,        --           .channel
			src6_startofpacket  => cmd_xbar_demux_src6_startofpacket,  --           .startofpacket
			src6_endofpacket    => cmd_xbar_demux_src6_endofpacket,    --           .endofpacket
			src7_ready          => cmd_xbar_demux_src7_ready,          --       src7.ready
			src7_valid          => cmd_xbar_demux_src7_valid,          --           .valid
			src7_data           => cmd_xbar_demux_src7_data,           --           .data
			src7_channel        => cmd_xbar_demux_src7_channel,        --           .channel
			src7_startofpacket  => cmd_xbar_demux_src7_startofpacket,  --           .startofpacket
			src7_endofpacket    => cmd_xbar_demux_src7_endofpacket,    --           .endofpacket
			src8_ready          => cmd_xbar_demux_src8_ready,          --       src8.ready
			src8_valid          => cmd_xbar_demux_src8_valid,          --           .valid
			src8_data           => cmd_xbar_demux_src8_data,           --           .data
			src8_channel        => cmd_xbar_demux_src8_channel,        --           .channel
			src8_startofpacket  => cmd_xbar_demux_src8_startofpacket,  --           .startofpacket
			src8_endofpacket    => cmd_xbar_demux_src8_endofpacket,    --           .endofpacket
			src9_ready          => cmd_xbar_demux_src9_ready,          --       src9.ready
			src9_valid          => cmd_xbar_demux_src9_valid,          --           .valid
			src9_data           => cmd_xbar_demux_src9_data,           --           .data
			src9_channel        => cmd_xbar_demux_src9_channel,        --           .channel
			src9_startofpacket  => cmd_xbar_demux_src9_startofpacket,  --           .startofpacket
			src9_endofpacket    => cmd_xbar_demux_src9_endofpacket,    --           .endofpacket
			src10_ready         => cmd_xbar_demux_src10_ready,         --      src10.ready
			src10_valid         => cmd_xbar_demux_src10_valid,         --           .valid
			src10_data          => cmd_xbar_demux_src10_data,          --           .data
			src10_channel       => cmd_xbar_demux_src10_channel,       --           .channel
			src10_startofpacket => cmd_xbar_demux_src10_startofpacket, --           .startofpacket
			src10_endofpacket   => cmd_xbar_demux_src10_endofpacket,   --           .endofpacket
			src11_ready         => cmd_xbar_demux_src11_ready,         --      src11.ready
			src11_valid         => cmd_xbar_demux_src11_valid,         --           .valid
			src11_data          => cmd_xbar_demux_src11_data,          --           .data
			src11_channel       => cmd_xbar_demux_src11_channel,       --           .channel
			src11_startofpacket => cmd_xbar_demux_src11_startofpacket, --           .startofpacket
			src11_endofpacket   => cmd_xbar_demux_src11_endofpacket,   --           .endofpacket
			src12_ready         => cmd_xbar_demux_src12_ready,         --      src12.ready
			src12_valid         => cmd_xbar_demux_src12_valid,         --           .valid
			src12_data          => cmd_xbar_demux_src12_data,          --           .data
			src12_channel       => cmd_xbar_demux_src12_channel,       --           .channel
			src12_startofpacket => cmd_xbar_demux_src12_startofpacket, --           .startofpacket
			src12_endofpacket   => cmd_xbar_demux_src12_endofpacket,   --           .endofpacket
			src13_ready         => cmd_xbar_demux_src13_ready,         --      src13.ready
			src13_valid         => cmd_xbar_demux_src13_valid,         --           .valid
			src13_data          => cmd_xbar_demux_src13_data,          --           .data
			src13_channel       => cmd_xbar_demux_src13_channel,       --           .channel
			src13_startofpacket => cmd_xbar_demux_src13_startofpacket, --           .startofpacket
			src13_endofpacket   => cmd_xbar_demux_src13_endofpacket,   --           .endofpacket
			src14_ready         => cmd_xbar_demux_src14_ready,         --      src14.ready
			src14_valid         => cmd_xbar_demux_src14_valid,         --           .valid
			src14_data          => cmd_xbar_demux_src14_data,          --           .data
			src14_channel       => cmd_xbar_demux_src14_channel,       --           .channel
			src14_startofpacket => cmd_xbar_demux_src14_startofpacket, --           .startofpacket
			src14_endofpacket   => cmd_xbar_demux_src14_endofpacket,   --           .endofpacket
			src15_ready         => cmd_xbar_demux_src15_ready,         --      src15.ready
			src15_valid         => cmd_xbar_demux_src15_valid,         --           .valid
			src15_data          => cmd_xbar_demux_src15_data,          --           .data
			src15_channel       => cmd_xbar_demux_src15_channel,       --           .channel
			src15_startofpacket => cmd_xbar_demux_src15_startofpacket, --           .startofpacket
			src15_endofpacket   => cmd_xbar_demux_src15_endofpacket,   --           .endofpacket
			src16_ready         => cmd_xbar_demux_src16_ready,         --      src16.ready
			src16_valid         => cmd_xbar_demux_src16_valid,         --           .valid
			src16_data          => cmd_xbar_demux_src16_data,          --           .data
			src16_channel       => cmd_xbar_demux_src16_channel,       --           .channel
			src16_startofpacket => cmd_xbar_demux_src16_startofpacket, --           .startofpacket
			src16_endofpacket   => cmd_xbar_demux_src16_endofpacket,   --           .endofpacket
			src17_ready         => cmd_xbar_demux_src17_ready,         --      src17.ready
			src17_valid         => cmd_xbar_demux_src17_valid,         --           .valid
			src17_data          => cmd_xbar_demux_src17_data,          --           .data
			src17_channel       => cmd_xbar_demux_src17_channel,       --           .channel
			src17_startofpacket => cmd_xbar_demux_src17_startofpacket, --           .startofpacket
			src17_endofpacket   => cmd_xbar_demux_src17_endofpacket,   --           .endofpacket
			src18_ready         => cmd_xbar_demux_src18_ready,         --      src18.ready
			src18_valid         => cmd_xbar_demux_src18_valid,         --           .valid
			src18_data          => cmd_xbar_demux_src18_data,          --           .data
			src18_channel       => cmd_xbar_demux_src18_channel,       --           .channel
			src18_startofpacket => cmd_xbar_demux_src18_startofpacket, --           .startofpacket
			src18_endofpacket   => cmd_xbar_demux_src18_endofpacket,   --           .endofpacket
			src19_ready         => cmd_xbar_demux_src19_ready,         --      src19.ready
			src19_valid         => cmd_xbar_demux_src19_valid,         --           .valid
			src19_data          => cmd_xbar_demux_src19_data,          --           .data
			src19_channel       => cmd_xbar_demux_src19_channel,       --           .channel
			src19_startofpacket => cmd_xbar_demux_src19_startofpacket, --           .startofpacket
			src19_endofpacket   => cmd_xbar_demux_src19_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_001 : component nios_ii_cmd_xbar_demux_001
		port map (
			clk                 => clk_100_clk,                            --        clk.clk
			reset               => rst_controller_reset_out_reset,         --  clk_reset.reset
			sink_ready          => limiter_001_cmd_src_ready,              --       sink.ready
			sink_channel        => limiter_001_cmd_src_channel,            --           .channel
			sink_data           => limiter_001_cmd_src_data,               --           .data
			sink_startofpacket  => limiter_001_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket    => limiter_001_cmd_src_endofpacket,        --           .endofpacket
			sink_valid          => limiter_001_cmd_valid_data,             -- sink_valid.data
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --       src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --           .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --           .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --           .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --           .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --           .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --       src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --           .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --           .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --           .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --           .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --           .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --       src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --           .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --           .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --           .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --           .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --           .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --       src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --           .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --           .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --           .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --           .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --           .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --       src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --           .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --           .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --           .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --           .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --           .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --       src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --           .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --           .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --           .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --           .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --           .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --       src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --           .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --           .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --           .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --           .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --           .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --       src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --           .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --           .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --           .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --           .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --           .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --       src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --           .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --           .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --           .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --           .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --           .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --       src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --           .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --           .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --           .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --           .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --           .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --      src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --           .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --           .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --           .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --           .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket,   --           .endofpacket
			src11_ready         => cmd_xbar_demux_001_src11_ready,         --      src11.ready
			src11_valid         => cmd_xbar_demux_001_src11_valid,         --           .valid
			src11_data          => cmd_xbar_demux_001_src11_data,          --           .data
			src11_channel       => cmd_xbar_demux_001_src11_channel,       --           .channel
			src11_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --           .startofpacket
			src11_endofpacket   => cmd_xbar_demux_001_src11_endofpacket,   --           .endofpacket
			src12_ready         => cmd_xbar_demux_001_src12_ready,         --      src12.ready
			src12_valid         => cmd_xbar_demux_001_src12_valid,         --           .valid
			src12_data          => cmd_xbar_demux_001_src12_data,          --           .data
			src12_channel       => cmd_xbar_demux_001_src12_channel,       --           .channel
			src12_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --           .startofpacket
			src12_endofpacket   => cmd_xbar_demux_001_src12_endofpacket,   --           .endofpacket
			src13_ready         => cmd_xbar_demux_001_src13_ready,         --      src13.ready
			src13_valid         => cmd_xbar_demux_001_src13_valid,         --           .valid
			src13_data          => cmd_xbar_demux_001_src13_data,          --           .data
			src13_channel       => cmd_xbar_demux_001_src13_channel,       --           .channel
			src13_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --           .startofpacket
			src13_endofpacket   => cmd_xbar_demux_001_src13_endofpacket,   --           .endofpacket
			src14_ready         => cmd_xbar_demux_001_src14_ready,         --      src14.ready
			src14_valid         => cmd_xbar_demux_001_src14_valid,         --           .valid
			src14_data          => cmd_xbar_demux_001_src14_data,          --           .data
			src14_channel       => cmd_xbar_demux_001_src14_channel,       --           .channel
			src14_startofpacket => cmd_xbar_demux_001_src14_startofpacket, --           .startofpacket
			src14_endofpacket   => cmd_xbar_demux_001_src14_endofpacket,   --           .endofpacket
			src15_ready         => cmd_xbar_demux_001_src15_ready,         --      src15.ready
			src15_valid         => cmd_xbar_demux_001_src15_valid,         --           .valid
			src15_data          => cmd_xbar_demux_001_src15_data,          --           .data
			src15_channel       => cmd_xbar_demux_001_src15_channel,       --           .channel
			src15_startofpacket => cmd_xbar_demux_001_src15_startofpacket, --           .startofpacket
			src15_endofpacket   => cmd_xbar_demux_001_src15_endofpacket,   --           .endofpacket
			src16_ready         => cmd_xbar_demux_001_src16_ready,         --      src16.ready
			src16_valid         => cmd_xbar_demux_001_src16_valid,         --           .valid
			src16_data          => cmd_xbar_demux_001_src16_data,          --           .data
			src16_channel       => cmd_xbar_demux_001_src16_channel,       --           .channel
			src16_startofpacket => cmd_xbar_demux_001_src16_startofpacket, --           .startofpacket
			src16_endofpacket   => cmd_xbar_demux_001_src16_endofpacket,   --           .endofpacket
			src17_ready         => cmd_xbar_demux_001_src17_ready,         --      src17.ready
			src17_valid         => cmd_xbar_demux_001_src17_valid,         --           .valid
			src17_data          => cmd_xbar_demux_001_src17_data,          --           .data
			src17_channel       => cmd_xbar_demux_001_src17_channel,       --           .channel
			src17_startofpacket => cmd_xbar_demux_001_src17_startofpacket, --           .startofpacket
			src17_endofpacket   => cmd_xbar_demux_001_src17_endofpacket,   --           .endofpacket
			src18_ready         => cmd_xbar_demux_001_src18_ready,         --      src18.ready
			src18_valid         => cmd_xbar_demux_001_src18_valid,         --           .valid
			src18_data          => cmd_xbar_demux_001_src18_data,          --           .data
			src18_channel       => cmd_xbar_demux_001_src18_channel,       --           .channel
			src18_startofpacket => cmd_xbar_demux_001_src18_startofpacket, --           .startofpacket
			src18_endofpacket   => cmd_xbar_demux_001_src18_endofpacket,   --           .endofpacket
			src19_ready         => cmd_xbar_demux_001_src19_ready,         --      src19.ready
			src19_valid         => cmd_xbar_demux_001_src19_valid,         --           .valid
			src19_data          => cmd_xbar_demux_001_src19_data,          --           .data
			src19_channel       => cmd_xbar_demux_001_src19_channel,       --           .channel
			src19_startofpacket => cmd_xbar_demux_001_src19_startofpacket, --           .startofpacket
			src19_endofpacket   => cmd_xbar_demux_001_src19_endofpacket,   --           .endofpacket
			src20_ready         => cmd_xbar_demux_001_src20_ready,         --      src20.ready
			src20_valid         => cmd_xbar_demux_001_src20_valid,         --           .valid
			src20_data          => cmd_xbar_demux_001_src20_data,          --           .data
			src20_channel       => cmd_xbar_demux_001_src20_channel,       --           .channel
			src20_startofpacket => cmd_xbar_demux_001_src20_startofpacket, --           .startofpacket
			src20_endofpacket   => cmd_xbar_demux_001_src20_endofpacket,   --           .endofpacket
			src21_ready         => cmd_xbar_demux_001_src21_ready,         --      src21.ready
			src21_valid         => cmd_xbar_demux_001_src21_valid,         --           .valid
			src21_data          => cmd_xbar_demux_001_src21_data,          --           .data
			src21_channel       => cmd_xbar_demux_001_src21_channel,       --           .channel
			src21_startofpacket => cmd_xbar_demux_001_src21_startofpacket, --           .startofpacket
			src21_endofpacket   => cmd_xbar_demux_001_src21_endofpacket,   --           .endofpacket
			src22_ready         => cmd_xbar_demux_001_src22_ready,         --      src22.ready
			src22_valid         => cmd_xbar_demux_001_src22_valid,         --           .valid
			src22_data          => cmd_xbar_demux_001_src22_data,          --           .data
			src22_channel       => cmd_xbar_demux_001_src22_channel,       --           .channel
			src22_startofpacket => cmd_xbar_demux_001_src22_startofpacket, --           .startofpacket
			src22_endofpacket   => cmd_xbar_demux_001_src22_endofpacket    --           .endofpacket
		);

	cmd_xbar_mux : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src3_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src3_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_004_src_data,             --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src4_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src4_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src4_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src4_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src4_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src4_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src4_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src4_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src4_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_005 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_005_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_005_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_005_src_data,             --          .data
			src_channel         => cmd_xbar_mux_005_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_005_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_005_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src5_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src5_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src5_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src5_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src5_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src5_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src5_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src5_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src5_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src5_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src5_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src5_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_006 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_006_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_006_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_006_src_data,             --          .data
			src_channel         => cmd_xbar_mux_006_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_006_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_006_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src6_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src6_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src6_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src6_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src6_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src6_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src6_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src6_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src6_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src6_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src6_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src6_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_007 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_007_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_007_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_007_src_data,             --          .data
			src_channel         => cmd_xbar_mux_007_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_007_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_007_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src7_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src7_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src7_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src7_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src7_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src7_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src7_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src7_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src7_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src7_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src7_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src7_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_008 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_008_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_008_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_008_src_data,             --          .data
			src_channel         => cmd_xbar_mux_008_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_008_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_008_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src8_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src8_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src8_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src8_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src8_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src8_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src8_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src8_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src8_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src8_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src8_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src8_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_009 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                           --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_009_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_009_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_009_src_data,             --          .data
			src_channel         => cmd_xbar_mux_009_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_009_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_009_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src9_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src9_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src9_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src9_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src9_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src9_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src9_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src9_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src9_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src9_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src9_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src9_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_010 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_010_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_010_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_010_src_data,              --          .data
			src_channel         => cmd_xbar_mux_010_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_010_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_010_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src10_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src10_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src10_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src10_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src10_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src10_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src10_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src10_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src10_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src10_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src10_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_011 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_011_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_011_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_011_src_data,              --          .data
			src_channel         => cmd_xbar_mux_011_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_011_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_011_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src11_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src11_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src11_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src11_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src11_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src11_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src11_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src11_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src11_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src11_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src11_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_012 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_012_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_012_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_012_src_data,              --          .data
			src_channel         => cmd_xbar_mux_012_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_012_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_012_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src12_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src12_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src12_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src12_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src12_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src12_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src12_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src12_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src12_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src12_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src12_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_013 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_013_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_013_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_013_src_data,              --          .data
			src_channel         => cmd_xbar_mux_013_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_013_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_013_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src13_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src13_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src13_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src13_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src13_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src13_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src13_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src13_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src13_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src13_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src13_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_014 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_014_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_014_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_014_src_data,              --          .data
			src_channel         => cmd_xbar_mux_014_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_014_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_014_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src14_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src14_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src14_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src14_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src14_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src14_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src14_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src14_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src14_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src14_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src14_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src14_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_015 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_015_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_015_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_015_src_data,              --          .data
			src_channel         => cmd_xbar_mux_015_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_015_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_015_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src15_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src15_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src15_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src15_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src15_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src15_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src15_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src15_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src15_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src15_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src15_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src15_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_016 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_016_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_016_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_016_src_data,              --          .data
			src_channel         => cmd_xbar_mux_016_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_016_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_016_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src16_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src16_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src16_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src16_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src16_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src16_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src16_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src16_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src16_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src16_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src16_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src16_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_017 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_017_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_017_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_017_src_data,              --          .data
			src_channel         => cmd_xbar_mux_017_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_017_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_017_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src17_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src17_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src17_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src17_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src17_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src17_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src17_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src17_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src17_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src17_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src17_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src17_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_018 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_018_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_018_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_018_src_data,              --          .data
			src_channel         => cmd_xbar_mux_018_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_018_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_018_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src18_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src18_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src18_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src18_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src18_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src18_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src18_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src18_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src18_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src18_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src18_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src18_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_019 : component nios_ii_cmd_xbar_mux
		port map (
			clk                 => clk_100_clk,                            --       clk.clk
			reset               => rst_controller_reset_out_reset,         -- clk_reset.reset
			src_ready           => cmd_xbar_mux_019_src_ready,             --       src.ready
			src_valid           => cmd_xbar_mux_019_src_valid,             --          .valid
			src_data            => cmd_xbar_mux_019_src_data,              --          .data
			src_channel         => cmd_xbar_mux_019_src_channel,           --          .channel
			src_startofpacket   => cmd_xbar_mux_019_src_startofpacket,     --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_019_src_endofpacket,       --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src19_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src19_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src19_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src19_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src19_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src19_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src19_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src19_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src19_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src19_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src19_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src19_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                       --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_005_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_005_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_005_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_005_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_005_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_006_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_006_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_006_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_006_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_006_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_007_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_007_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_007_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_007_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_007_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_007_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_008_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_008_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_008_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_008_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_008_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_008_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_009_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_009_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_009_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_009_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_009_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_009_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_010_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_010_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_010_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_010_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_010_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_010_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_011_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_011_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_011_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_011_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_011_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_011_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_012_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_012_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_012_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_012_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_012_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_012_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_013_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_013_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_013_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_013_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_013_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_013_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_014_src_ready,               --      sink.ready
			sink_channel       => id_router_014_src_channel,             --          .channel
			sink_data          => id_router_014_src_data,                --          .data
			sink_startofpacket => id_router_014_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_014_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_014_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_014_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_014_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_014_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_014_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_014_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_014_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_015 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_015_src_ready,               --      sink.ready
			sink_channel       => id_router_015_src_channel,             --          .channel
			sink_data          => id_router_015_src_data,                --          .data
			sink_startofpacket => id_router_015_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_015_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_015_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_015_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_015_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_015_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_015_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_015_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_015_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_015_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_015_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_016 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_016_src_ready,               --      sink.ready
			sink_channel       => id_router_016_src_channel,             --          .channel
			sink_data          => id_router_016_src_data,                --          .data
			sink_startofpacket => id_router_016_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_016_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_016_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_016_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_016_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_016_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_016_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_016_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_016_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_016_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_016_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_016_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_017 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_017_src_ready,               --      sink.ready
			sink_channel       => id_router_017_src_channel,             --          .channel
			sink_data          => id_router_017_src_data,                --          .data
			sink_startofpacket => id_router_017_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_017_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_017_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_017_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_017_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_017_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_017_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_017_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_017_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_017_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_017_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_017_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_018 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_018_src_ready,               --      sink.ready
			sink_channel       => id_router_018_src_channel,             --          .channel
			sink_data          => id_router_018_src_data,                --          .data
			sink_startofpacket => id_router_018_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_018_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_018_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_018_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_018_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_018_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_018_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_018_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_018_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_018_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_018_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_018_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_018_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_018_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_018_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_019 : component nios_ii_rsp_xbar_demux
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_019_src_ready,               --      sink.ready
			sink_channel       => id_router_019_src_channel,             --          .channel
			sink_data          => id_router_019_src_data,                --          .data
			sink_startofpacket => id_router_019_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_019_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_019_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_019_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_019_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_019_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_019_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_019_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_019_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_019_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_019_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_019_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_019_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_019_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_019_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_020 : component nios_ii_rsp_xbar_demux_020
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_020_src_ready,               --      sink.ready
			sink_channel       => id_router_020_src_channel,             --          .channel
			sink_data          => id_router_020_src_data,                --          .data
			sink_startofpacket => id_router_020_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_020_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_020_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_020_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_020_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_020_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_020_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_020_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_020_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_021 : component nios_ii_rsp_xbar_demux_020
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_003_src_ready,           --      sink.ready
			sink_channel       => width_adapter_003_src_channel,         --          .channel
			sink_data          => width_adapter_003_src_data,            --          .data
			sink_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_003_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_021_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_021_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_021_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_021_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_021_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_021_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_022 : component nios_ii_rsp_xbar_demux_020
		port map (
			clk                => clk_100_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_022_src_ready,               --      sink.ready
			sink_channel       => id_router_022_src_channel,             --          .channel
			sink_data          => id_router_022_src_data,                --          .data
			sink_startofpacket => id_router_022_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_022_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_022_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_022_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_022_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_022_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_022_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_022_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_022_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component nios_ii_rsp_xbar_mux
		port map (
			clk                  => clk_100_clk,                           --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid            => rsp_xbar_mux_src_valid,                --          .valid
			src_data             => rsp_xbar_mux_src_data,                 --          .data
			src_channel          => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket    => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink14_ready         => rsp_xbar_demux_014_src0_ready,         --    sink14.ready
			sink14_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink14_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink14_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink14_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink14_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			sink15_ready         => rsp_xbar_demux_015_src0_ready,         --    sink15.ready
			sink15_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			sink15_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			sink15_data          => rsp_xbar_demux_015_src0_data,          --          .data
			sink15_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			sink15_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			sink16_ready         => rsp_xbar_demux_016_src0_ready,         --    sink16.ready
			sink16_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			sink16_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			sink16_data          => rsp_xbar_demux_016_src0_data,          --          .data
			sink16_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			sink16_endofpacket   => rsp_xbar_demux_016_src0_endofpacket,   --          .endofpacket
			sink17_ready         => rsp_xbar_demux_017_src0_ready,         --    sink17.ready
			sink17_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			sink17_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			sink17_data          => rsp_xbar_demux_017_src0_data,          --          .data
			sink17_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			sink17_endofpacket   => rsp_xbar_demux_017_src0_endofpacket,   --          .endofpacket
			sink18_ready         => rsp_xbar_demux_018_src0_ready,         --    sink18.ready
			sink18_valid         => rsp_xbar_demux_018_src0_valid,         --          .valid
			sink18_channel       => rsp_xbar_demux_018_src0_channel,       --          .channel
			sink18_data          => rsp_xbar_demux_018_src0_data,          --          .data
			sink18_startofpacket => rsp_xbar_demux_018_src0_startofpacket, --          .startofpacket
			sink18_endofpacket   => rsp_xbar_demux_018_src0_endofpacket,   --          .endofpacket
			sink19_ready         => rsp_xbar_demux_019_src0_ready,         --    sink19.ready
			sink19_valid         => rsp_xbar_demux_019_src0_valid,         --          .valid
			sink19_channel       => rsp_xbar_demux_019_src0_channel,       --          .channel
			sink19_data          => rsp_xbar_demux_019_src0_data,          --          .data
			sink19_startofpacket => rsp_xbar_demux_019_src0_startofpacket, --          .startofpacket
			sink19_endofpacket   => rsp_xbar_demux_019_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component nios_ii_rsp_xbar_mux_001
		port map (
			clk                  => clk_100_clk,                           --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src1_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src1_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src1_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src1_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src1_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src1_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src1_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src1_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src1_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src1_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src1_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src1_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src1_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src1_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src1_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src1_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src1_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src1_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src1_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src1_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src1_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src1_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src1_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src1_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src1_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src1_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src1_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src1_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src1_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src1_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src1_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src1_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src1_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src1_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src1_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src1_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src1_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src1_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src1_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src1_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src1_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src1_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src1_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src1_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src1_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src1_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src1_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src1_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src1_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src1_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src1_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src1_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src1_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src1_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src1_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src1_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src1_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src1_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src1_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src1_endofpacket,   --          .endofpacket
			sink14_ready         => rsp_xbar_demux_014_src1_ready,         --    sink14.ready
			sink14_valid         => rsp_xbar_demux_014_src1_valid,         --          .valid
			sink14_channel       => rsp_xbar_demux_014_src1_channel,       --          .channel
			sink14_data          => rsp_xbar_demux_014_src1_data,          --          .data
			sink14_startofpacket => rsp_xbar_demux_014_src1_startofpacket, --          .startofpacket
			sink14_endofpacket   => rsp_xbar_demux_014_src1_endofpacket,   --          .endofpacket
			sink15_ready         => rsp_xbar_demux_015_src1_ready,         --    sink15.ready
			sink15_valid         => rsp_xbar_demux_015_src1_valid,         --          .valid
			sink15_channel       => rsp_xbar_demux_015_src1_channel,       --          .channel
			sink15_data          => rsp_xbar_demux_015_src1_data,          --          .data
			sink15_startofpacket => rsp_xbar_demux_015_src1_startofpacket, --          .startofpacket
			sink15_endofpacket   => rsp_xbar_demux_015_src1_endofpacket,   --          .endofpacket
			sink16_ready         => rsp_xbar_demux_016_src1_ready,         --    sink16.ready
			sink16_valid         => rsp_xbar_demux_016_src1_valid,         --          .valid
			sink16_channel       => rsp_xbar_demux_016_src1_channel,       --          .channel
			sink16_data          => rsp_xbar_demux_016_src1_data,          --          .data
			sink16_startofpacket => rsp_xbar_demux_016_src1_startofpacket, --          .startofpacket
			sink16_endofpacket   => rsp_xbar_demux_016_src1_endofpacket,   --          .endofpacket
			sink17_ready         => rsp_xbar_demux_017_src1_ready,         --    sink17.ready
			sink17_valid         => rsp_xbar_demux_017_src1_valid,         --          .valid
			sink17_channel       => rsp_xbar_demux_017_src1_channel,       --          .channel
			sink17_data          => rsp_xbar_demux_017_src1_data,          --          .data
			sink17_startofpacket => rsp_xbar_demux_017_src1_startofpacket, --          .startofpacket
			sink17_endofpacket   => rsp_xbar_demux_017_src1_endofpacket,   --          .endofpacket
			sink18_ready         => rsp_xbar_demux_018_src1_ready,         --    sink18.ready
			sink18_valid         => rsp_xbar_demux_018_src1_valid,         --          .valid
			sink18_channel       => rsp_xbar_demux_018_src1_channel,       --          .channel
			sink18_data          => rsp_xbar_demux_018_src1_data,          --          .data
			sink18_startofpacket => rsp_xbar_demux_018_src1_startofpacket, --          .startofpacket
			sink18_endofpacket   => rsp_xbar_demux_018_src1_endofpacket,   --          .endofpacket
			sink19_ready         => rsp_xbar_demux_019_src1_ready,         --    sink19.ready
			sink19_valid         => rsp_xbar_demux_019_src1_valid,         --          .valid
			sink19_channel       => rsp_xbar_demux_019_src1_channel,       --          .channel
			sink19_data          => rsp_xbar_demux_019_src1_data,          --          .data
			sink19_startofpacket => rsp_xbar_demux_019_src1_startofpacket, --          .startofpacket
			sink19_endofpacket   => rsp_xbar_demux_019_src1_endofpacket,   --          .endofpacket
			sink20_ready         => rsp_xbar_demux_020_src0_ready,         --    sink20.ready
			sink20_valid         => rsp_xbar_demux_020_src0_valid,         --          .valid
			sink20_channel       => rsp_xbar_demux_020_src0_channel,       --          .channel
			sink20_data          => rsp_xbar_demux_020_src0_data,          --          .data
			sink20_startofpacket => rsp_xbar_demux_020_src0_startofpacket, --          .startofpacket
			sink20_endofpacket   => rsp_xbar_demux_020_src0_endofpacket,   --          .endofpacket
			sink21_ready         => rsp_xbar_demux_021_src0_ready,         --    sink21.ready
			sink21_valid         => rsp_xbar_demux_021_src0_valid,         --          .valid
			sink21_channel       => rsp_xbar_demux_021_src0_channel,       --          .channel
			sink21_data          => rsp_xbar_demux_021_src0_data,          --          .data
			sink21_startofpacket => rsp_xbar_demux_021_src0_startofpacket, --          .startofpacket
			sink21_endofpacket   => rsp_xbar_demux_021_src0_endofpacket,   --          .endofpacket
			sink22_ready         => rsp_xbar_demux_022_src0_ready,         --    sink22.ready
			sink22_valid         => rsp_xbar_demux_022_src0_valid,         --          .valid
			sink22_channel       => rsp_xbar_demux_022_src0_channel,       --          .channel
			sink22_data          => rsp_xbar_demux_022_src0_data,          --          .data
			sink22_startofpacket => rsp_xbar_demux_022_src0_startofpacket, --          .startofpacket
			sink22_endofpacket   => rsp_xbar_demux_022_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component nios_ii_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 56,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 65,
			IN_PKT_BYTE_CNT_L             => 63,
			IN_PKT_TRANS_COMPRESSED_READ  => 57,
			IN_PKT_BURSTWRAP_H            => 68,
			IN_PKT_BURSTWRAP_L            => 66,
			IN_PKT_BURST_SIZE_H           => 71,
			IN_PKT_BURST_SIZE_L           => 69,
			IN_PKT_RESPONSE_STATUS_H      => 97,
			IN_PKT_RESPONSE_STATUS_L      => 96,
			IN_PKT_TRANS_EXCLUSIVE        => 62,
			IN_PKT_BURST_TYPE_H           => 73,
			IN_PKT_BURST_TYPE_L           => 72,
			IN_ST_DATA_W                  => 98,
			OUT_PKT_ADDR_H                => 38,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 47,
			OUT_PKT_BYTE_CNT_L            => 45,
			OUT_PKT_TRANS_COMPRESSED_READ => 39,
			OUT_PKT_BURST_SIZE_H          => 53,
			OUT_PKT_BURST_SIZE_L          => 51,
			OUT_PKT_RESPONSE_STATUS_H     => 79,
			OUT_PKT_RESPONSE_STATUS_L     => 78,
			OUT_PKT_TRANS_EXCLUSIVE       => 44,
			OUT_PKT_BURST_TYPE_H          => 55,
			OUT_PKT_BURST_TYPE_L          => 54,
			OUT_ST_DATA_W                 => 80,
			ST_CHANNEL_W                  => 23,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_100_clk,                        --       clk.clk
			reset                => rst_controller_reset_out_reset,     -- clk_reset.reset
			in_valid             => cmd_xbar_mux_001_src_valid,         --      sink.valid
			in_channel           => cmd_xbar_mux_001_src_channel,       --          .channel
			in_startofpacket     => cmd_xbar_mux_001_src_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_001_src_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_mux_001_src_ready,         --          .ready
			in_data              => cmd_xbar_mux_001_src_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component nios_ii_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 38,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 47,
			IN_PKT_BYTE_CNT_L             => 45,
			IN_PKT_TRANS_COMPRESSED_READ  => 39,
			IN_PKT_BURSTWRAP_H            => 50,
			IN_PKT_BURSTWRAP_L            => 48,
			IN_PKT_BURST_SIZE_H           => 53,
			IN_PKT_BURST_SIZE_L           => 51,
			IN_PKT_RESPONSE_STATUS_H      => 79,
			IN_PKT_RESPONSE_STATUS_L      => 78,
			IN_PKT_TRANS_EXCLUSIVE        => 44,
			IN_PKT_BURST_TYPE_H           => 55,
			IN_PKT_BURST_TYPE_L           => 54,
			IN_ST_DATA_W                  => 80,
			OUT_PKT_ADDR_H                => 56,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 65,
			OUT_PKT_BYTE_CNT_L            => 63,
			OUT_PKT_TRANS_COMPRESSED_READ => 57,
			OUT_PKT_BURST_SIZE_H          => 71,
			OUT_PKT_BURST_SIZE_L          => 69,
			OUT_PKT_RESPONSE_STATUS_H     => 97,
			OUT_PKT_RESPONSE_STATUS_L     => 96,
			OUT_PKT_TRANS_EXCLUSIVE       => 62,
			OUT_PKT_BURST_TYPE_H          => 73,
			OUT_PKT_BURST_TYPE_L          => 72,
			OUT_ST_DATA_W                 => 98,
			ST_CHANNEL_W                  => 23,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_100_clk,                         --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_001_src_valid,             --      sink.valid
			in_channel           => id_router_001_src_channel,           --          .channel
			in_startofpacket     => id_router_001_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_001_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_001_src_ready,             --          .ready
			in_data              => id_router_001_src_data,              --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_002 : component nios_ii_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 56,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 65,
			IN_PKT_BYTE_CNT_L             => 63,
			IN_PKT_TRANS_COMPRESSED_READ  => 57,
			IN_PKT_BURSTWRAP_H            => 68,
			IN_PKT_BURSTWRAP_L            => 66,
			IN_PKT_BURST_SIZE_H           => 71,
			IN_PKT_BURST_SIZE_L           => 69,
			IN_PKT_RESPONSE_STATUS_H      => 97,
			IN_PKT_RESPONSE_STATUS_L      => 96,
			IN_PKT_TRANS_EXCLUSIVE        => 62,
			IN_PKT_BURST_TYPE_H           => 73,
			IN_PKT_BURST_TYPE_L           => 72,
			IN_ST_DATA_W                  => 98,
			OUT_PKT_ADDR_H                => 38,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 47,
			OUT_PKT_BYTE_CNT_L            => 45,
			OUT_PKT_TRANS_COMPRESSED_READ => 39,
			OUT_PKT_BURST_SIZE_H          => 53,
			OUT_PKT_BURST_SIZE_L          => 51,
			OUT_PKT_RESPONSE_STATUS_H     => 79,
			OUT_PKT_RESPONSE_STATUS_L     => 78,
			OUT_PKT_TRANS_EXCLUSIVE       => 44,
			OUT_PKT_BURST_TYPE_H          => 55,
			OUT_PKT_BURST_TYPE_L          => 54,
			OUT_ST_DATA_W                 => 80,
			ST_CHANNEL_W                  => 23,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_100_clk,                            --       clk.clk
			reset                => rst_controller_reset_out_reset,         -- clk_reset.reset
			in_valid             => cmd_xbar_demux_001_src21_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_001_src21_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_001_src21_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_001_src21_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_001_src21_ready,         --          .ready
			in_data              => cmd_xbar_demux_001_src21_data,          --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_002_src_data,             --          .data
			out_channel          => width_adapter_002_src_channel,          --          .channel
			out_valid            => width_adapter_002_src_valid,            --          .valid
			out_ready            => width_adapter_002_src_ready,            --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                                   -- (terminated)
		);

	width_adapter_003 : component nios_ii_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 38,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 47,
			IN_PKT_BYTE_CNT_L             => 45,
			IN_PKT_TRANS_COMPRESSED_READ  => 39,
			IN_PKT_BURSTWRAP_H            => 50,
			IN_PKT_BURSTWRAP_L            => 48,
			IN_PKT_BURST_SIZE_H           => 53,
			IN_PKT_BURST_SIZE_L           => 51,
			IN_PKT_RESPONSE_STATUS_H      => 79,
			IN_PKT_RESPONSE_STATUS_L      => 78,
			IN_PKT_TRANS_EXCLUSIVE        => 44,
			IN_PKT_BURST_TYPE_H           => 55,
			IN_PKT_BURST_TYPE_L           => 54,
			IN_ST_DATA_W                  => 80,
			OUT_PKT_ADDR_H                => 56,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 65,
			OUT_PKT_BYTE_CNT_L            => 63,
			OUT_PKT_TRANS_COMPRESSED_READ => 57,
			OUT_PKT_BURST_SIZE_H          => 71,
			OUT_PKT_BURST_SIZE_L          => 69,
			OUT_PKT_RESPONSE_STATUS_H     => 97,
			OUT_PKT_RESPONSE_STATUS_L     => 96,
			OUT_PKT_TRANS_EXCLUSIVE       => 62,
			OUT_PKT_BURST_TYPE_H          => 73,
			OUT_PKT_BURST_TYPE_L          => 72,
			OUT_ST_DATA_W                 => 98,
			ST_CHANNEL_W                  => 23,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_100_clk,                         --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_021_src_valid,             --      sink.valid
			in_channel           => id_router_021_src_channel,           --          .channel
			in_startofpacket     => id_router_021_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_021_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_021_src_ready,             --          .ready
			in_data              => id_router_021_src_data,              --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_003_src_data,          --          .data
			out_channel          => width_adapter_003_src_channel,       --          .channel
			out_valid            => width_adapter_003_src_valid,         --          .valid
			out_ready            => width_adapter_003_src_ready,         --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	irq_mapper : component nios_ii_irq_mapper
		port map (
			clk           => clk_100_clk,                    --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,       -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_irq,       -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_irq,       -- receiver7.irq
			receiver8_irq => irq_mapper_receiver8_irq,       -- receiver8.irq
			sender_irq    => nios2_qsys_0_d_irq_irq          --    sender.irq
		);

	reset_100_reset_n_ports_inv <= not reset_100_reset_n;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	audio_sos_s1_translator_avalon_anti_slave_0_write_ports_inv <= not audio_sos_s1_translator_avalon_anti_slave_0_write;

	dac_irq_s1_translator_avalon_anti_slave_0_write_ports_inv <= not dac_irq_s1_translator_avalon_anti_slave_0_write;

	clap_irq_s1_translator_avalon_anti_slave_0_write_ports_inv <= not clap_irq_s1_translator_avalon_anti_slave_0_write;

	hh_irq_s1_translator_avalon_anti_slave_0_write_ports_inv <= not hh_irq_s1_translator_avalon_anti_slave_0_write;

	snare_irq_s1_translator_avalon_anti_slave_0_write_ports_inv <= not snare_irq_s1_translator_avalon_anti_slave_0_write;

	kick_irq_s1_translator_avalon_anti_slave_0_write_ports_inv <= not kick_irq_s1_translator_avalon_anti_slave_0_write;

	kb_irq_s1_translator_avalon_anti_slave_0_write_ports_inv <= not kb_irq_s1_translator_avalon_anti_slave_0_write;

	seq_hh_s1_translator_avalon_anti_slave_0_write_ports_inv <= not seq_hh_s1_translator_avalon_anti_slave_0_write;

	seq_snare_s1_translator_avalon_anti_slave_0_write_ports_inv <= not seq_snare_s1_translator_avalon_anti_slave_0_write;

	led_r_s1_translator_avalon_anti_slave_0_write_ports_inv <= not led_r_s1_translator_avalon_anti_slave_0_write;

	timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_0_s1_translator_avalon_anti_slave_0_write;

	seq_clap_s1_translator_avalon_anti_slave_0_write_ports_inv <= not seq_clap_s1_translator_avalon_anti_slave_0_write;

	seq_kick_s1_translator_avalon_anti_slave_0_write_ports_inv <= not seq_kick_s1_translator_avalon_anti_slave_0_write;

	wr_address_s1_translator_avalon_anti_slave_0_write_ports_inv <= not wr_address_s1_translator_avalon_anti_slave_0_write;

	color_out_s1_translator_avalon_anti_slave_0_write_ports_inv <= not color_out_s1_translator_avalon_anti_slave_0_write;

	wr_en_s1_translator_avalon_anti_slave_0_write_ports_inv <= not wr_en_s1_translator_avalon_anti_slave_0_write;

	timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_1_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of nios_ii
